`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
UTEFCZ1BkAWC+zJiq9ChFr4TKVPHHZn0ihyu1/CgZ3/SHXsfmegpf1MbYSz7xmhY
9h27mXjFutADvqE6m9JwjvR4jl7hx+j+kV2+7wJU3UQOv203MeuVYEGXTmdm/iaJ
OMmajbR26rMjk1L6RUxSHo9yAmM6OUut9nCN39yzKxg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 749632)
oTPQST9QdV3iOnHampCWrSm01LNwe2JPwYhF22RRTlSfoE8IMWYXhWIyPez8sRFz
4U5NCgUPrUqG/oYEW1EDN1EemUTF1m0d1U6J2juJzQy8h8f7GY82+EGBIo70POfX
KdNgmStdw+FiPwFf83NMNoAAmYz62Oravyj8rhoV4RQG6G9pJ3kfp5ZTsuft2PZs
hv9I9B9pDMwo7hVwRZQfLsk87OCUObUwg9Poyb1OeTvZ9NzjC8fphLAOiutBYrW9
sE1MtRWvBMe5cJCEH2qYHdAm3JPowai5Z7Yd55cE/NtJilGH4BLrxwbFyIbslqk/
l+47PEcBCUxuf5IW+k2HE4RSNTMi08G8HxnEMshtrbiOi1yMlI7adHS4NAF+NGy1
FXNdbahTiKUv9Ru58jtKzsoOg+PEKvQf0LbWqqIBW69zk+qroGo/h0DyMCxEfhsn
3eLC/9WvRkDV7SwnQFy0w7+DeKXK4vGhyqBb5urxrsiUtQ1pxKgEsj7kr3/AVWH1
iP3JaHKVOQthnPO1we8NTRSEC1hX3FV/sJ7fkUcEWWSOD3rAEA1n+zS4CriCXND3
M7VGc1BYEVVmJVR/w2PH/GeOkAWxZSOX39QKoGnGhGuUBKo6aw9Oz032AsvvIo/q
yoDVswqOtoVC4JchW1w4ENBz1w+6oyq13H3N3vHeglXnzFWhnWsKQ0DLnE+A30uP
8hlmOKAt1H5glko6y3ZQ/H+1Ct56O9mHRH5vh8MQ+pXYIEL5XFf4b9n0CYWb87qZ
wq61wrtfY5DXte4fVf6dYNtuBPhecjdL76E0GF1BKeUOWvh6CuyZIic/LvwAoGO1
YqRXDMFA0Q4+pISTSNBuzqfJb0rWbouiZIrjEJjGxM5gl63KXhBoe1RhgORoARbI
PtW+o0YJIchwMyvS4U42zx3zkEyc6/mKd+PkXM+P5hKa/Qdza2hpuCSN1HkKSNta
myVLO+V60XIKxi0x/t305RZeevNoURzwnQ8Qih4xY/BVyTK7VofolfStCkdvf3tA
K/+r3ilF7irVCo9JiDLIc6VDzshKnLi7Bys6jTEV9AFk1iTQUUNY7R/vmYVQWm2A
tgvjjcYPvzUDVx/B7R+tbgzt5EsR3BEOexCiE4bUjnxJZ0IK/DyUCUGvIUR5x9jP
v/w58I8eGTHygUqHb9qu6AqdwCOJGPsyEEcpcPAVtgS76kjwluvmj3W5BORlR8eQ
66cLQrne8ynXlxNrjAWANwqBqB8WuoUTS9Ulnl0Bg0wZEb9uua8pFJX8diIwOy6X
OVByMM6rdPaAWmNKozCqS2eG+KFs8qQtBE7Yz3hE/3D4eHfOTBu/vQv2Jxv2gyf4
Q1pIWpJepF/4ATzwK/3jnDHvPjJ42MTUtdsikzfK1n2VzZPms9ctJPw3yVfgR/Nq
0m5821XXxiGvMWjoCX3XuFBcmxgrOQ61dVmTlhtfl5SYup7vcZDpy4trYvqDOr/N
kBuDVIA/MOSBImIZl9pfhEYCtn9nZ8GIWziBODvZThyHiD8BQDixlZywhd55OZC5
zD+OeL/3qaSh1ULxQWOOz93yQK3e3oh3oMs1RYPSI0kw4NahZtbjsADC4nqq8fP3
NNHCnfXIKUdwcBa02pAm+FE+3/ZM1cwtU2bfBp7d6IwtJHkpa8mfPxT6Nyut79v/
tYE5EVHpIv2r7YBMeYE71aSPxGWK63uuoI0eJbim8GJtXm4MHKwpaOtS5zgGVlkF
2fCk0C+m1rk/c4exduuWk3Ffb+3+4IUS25RJeZepuqitXDojyv2edfka+afwWAp0
gxEsdskrQMuPovT6Yt5Rbe7CEHsguVtolDkVlYGM++v+AjlWOfEB4xdBrPUTffZa
sjS9y9Yb8LL/rCzk3tRB4mjCaaaL+Puv/WYRQ3TBvceY+VktWuKn96AsPzPl4Tin
WaRvq6XGlSP58bRbYR51BNjIjMlIxDGC612cScJJOJJPFRAU4h7KDU1q2NNAEjEC
SZb2n8as9fb0WrqyzBNPX7Ksy6PrMHPaOTfKfd5SyZWuCcq05GIrytlHOnQpsXc+
PP/Afh6rihQAOquaidw4C5DBCLMbKGMRrOBUTFQA3OKn/s0rnrBkuAdDvAFyzu0d
JsWkHu3nzSotrL6wWGC7+uOaEsXOt9ZqzVHriimJaAH/3daOhKtPlvo49F5EWty8
eY5GYA8I0df4P3xsQ/lhVsZzBuHa4qcuSVjdijcd0r2fiInu+uGpnzBjkD0fIudU
GW9q675LvuJVHY/xICTKSUQqos+Ub/hYzboJM8m9vOgnVUh7hnu2jGioQijCR1Sy
GKgtk1qrZuiPIOkBXrksjU9w8Ac/PoyreRf7pZFEjszgSWBVPlZ2RjheVbUKqTuT
VCzs4PMCxv2aOOvwcxUiP/7J2WoU3rMYGu1UkMD+CCkFKBw2Q816nIWk1mUvobH9
alhRs5sNoJUorE513M3EbnXloRH6/TkiDSORXPQURcQCjX+BJqMZgG3m4NbKQfQ5
R8BudLmedEdoQxwGKGnRHLATL/tSlKkg0ZwKQi9NMuAF9n6usaanFEi9pt65bO/P
B23o+JD4qAOQHY5kdfyV/B0tLuhk42toBM7eH3aqRONUivJL02XVSqmbH3qqN9dP
DLgtzd8reqjRScGnejR3By9bv18kPzA52NYY86xvstUH8/gyRJhW8dwTe4A64FNV
z2O4SleL9jFM/55J13PGq73H5Rfz6NYKFHK0pdONJNOLVp72BMttDWfUlWtQQjUI
/ZbjF0HgMnHBkdkMZAspTjcRbMcYD6psiHcgr4RCHXitt/74q2L2OYB064yyWIPX
8PpXtRSgbHvgSGzOhitZFd8nQUAAN00PN6lSQm1VldFqpOsdKDFLgwjw96TGN6d9
Pp4ustjm1e/eMRmqcYXYuSzOU2RcvY3f+jVWqKIp0ZW+udidIYn5blQGJUBzKqDz
TGSdIhj9rt23y9pvs7hIRcyl9ikDEy7IiVt3c9TfsSiVjNmYcSXpQIF0+s/TPL8P
D7tlqcvXICyav33dseu4gsSgQLmituck4DjKBVux010jz38FGUuf2XYKHt/aIcGG
iAHHbDsmx3YdGxVMZAB5un/3uPisEY4imH2uKgdg3Sut+adx9HxvfSTcZ8+o0qUt
9pH2QqvHch04RlYZdafegTYs8ryZTuIypFJYDo5v+tZSX25CMLRF1XUGThkiWWbd
7RBDmaWZhcW5lBdJ74EmOBOP3aXcVFma8MZdP7nK15KuC8ksN3tD83r0oE522xUd
JGCYCOGCvc/54TWEx3W3ELB5vq3KJ7Nq1AQGwKI1hpsq3U4eq6AxMPW6UmY+eEY7
vpB1zOC903Q6BT8nDHZlA6iMEYf0iJa9yzk+ghUTZYyK/poYrzxMaMOSliR449Z7
xpx9ki++D+gvkfsHFfPI3elfmKZe6QnQFSQaGaPk/xjHle2HpABSC7tdWKhy8xTS
3UPmGUQ7rywp27K+EBMhNCf0wwXNPcRNL5d9jTe7NEveKZ48TGYBxCZMRzevm0pC
THNkon69DSEA8BaYVIzElPJLK3POgbP+RqIhqaknJe5t65557ylzRzs6tbCcfh7D
gA1/25AZk5m9kbCVeDJ+2wJiHJGUfH3lqCibPVTi2bdwmECRNPOHtkhG7DS3wTy9
8nUAZJlyJlACEHr/e1od8wljouQI2aoqGJeaSqTCFW9v3/pqIWyzKeGzxZHIsJad
xDexCid/lRK37scrU5Qol0Cnud8r9uwvEe66B4Fizxn1pqCR9ETWbtSuCaDDWsRA
fx3uvabGARv0iVpfv8ns6+K/L9s+c8iS4jYWUlkUHe2Adkwvxb1zMkfNgayx4Pgy
+Mn1SvdjevyNVQqH6BNid1Oyvws0zvwp0lYUu7N1YL5bG83uGnRxauj3eoGr8JHd
t6eB8xNDi4335E1O/xpvBmjENj0WXAui/2v7E2aeZvFmy7vcffLoBC0GnYALu+3i
UTkgWWU5WBqKJHkUq0JUNWvVdHIXHIuO8txVBjL0MUNYVHI0lFdcantr4P/iFXrG
X3DbsnI9XsfcB42p7K12SwkqDIqpYgK7pfpK1gHIERK37dmUfEys1ifT10uXVYqZ
p/Zmk68FM8d3Bw8hwc6FG1NkKNrKlMIAv6aHjsVosbjuSpL+aDruT5GZG9k4Qhkz
lsgfmJob2aZea+ErZmnWoQ/04uvhd5hU6HdUC0QAcTyzsUCBBnjN03iHWNx51H+h
uMAXwckIvMOzdxMdP5duG9czBbhS+2M7VzVoGKb6r5GA+aBp6Ts6HEQuxeX/Y+Ri
WogDh7Uh9iD5O2g5Zs95TLL2wERGH/pHIA7QX31Bzj6xalOwfvvweU89IwH8gjZd
PfYUjiuWbkbwME74kaq/g/LT8HNxOI/QgOgeetHrfRyj3QU59+bFVqXqNPLuAdRL
Vn0siE5vjUSJGpMw/Ocf83AcHHt1805ri1/d0uvLjTgBOVDtEPONm8yyODfbiQzE
/joYkvpnzE5+ksErSq0XtRf7EqSQ6mBgEGwNtPTP9jepjt/8A7T+/RQ3pF0KKpyu
zS11O/FoN4JdR9pUIC7h0R5GaNxNkQ3X+QuaLGQGslf5yRAw5FCwjsQ8qGQHd26m
kMoEuDgpsqxFeONlKRuKbv/gnqneiPQ4FFKN6Ar4dbJgteOuWj7fIAnX9zWNHfic
xYvHh+126tUVzDxLrQ2WldhJbadST+SorF5y4rY1yHX8hyKXmhCESIdlEfIXR55Z
W2g++VLkcNglXO1/j9UU90vJcc/KAHxlhIJl6hYT6Jjk6fyHHMfu+qeItU6C2ivy
Q7kRGdT+o1STmt7GRL27I5Pmt6u8a1Dt3aTK5RpT495p9dnbdKrM3bKLExgr79OT
YM/+qu8M/5ke6qWstHyoj9UFTg217H72SxMZ4/C3rpdXaHuxSvuXOUILCJj0KNn9
6Lbv5AJBAB/8xTKBLv0H81yP1dTIFiDjm1WCycD5BkyDmHFKdSj9MsAivEODPSdp
Q+yCuBhJpkxSx63v6vMiRow0WorBkCwAIHNxfXLBdfycY/XjSAOERhjKiwBaN0bP
xptcrJbS3+CxfFms7cuT06Q70pUYWr+36HnC50IQlsfiYfOBCHzFWfnYXBkPLnBT
1afNxwPClp+LXA1zx1Kc6YI/5MSBacwsE4KH2Zq7BzfVuvFaBWqlRrxUowpnaeOX
1wJ1rIPETI9mmhVssedNLJX5K/RORYLwiq2SHmveQsQpwTlyEqVdSLDaiAcQ9gYs
AKfQv0iit0+sfcK47xb0o7UZwTQbA4Sl3qP2mM6LYtthcsXLVhBDuSaQXzcEc38y
aa1J7KHVM3KiMNNBtgDDZ7Bz229o+lNBj7nZ/vjdqQG86cMxf0b+wVFVWKWaWj3V
q0tZYqzL5SQ5f5aAV50IEbaFja9qZRsbjGnbOzWNEC3S4srzv4UhUAqpIgTNjS9l
48OUznwEdxDD5xyVmTgbaKhdn0fxsc687niyp0+vZ1dUfgd2jRZsdPVwklOd9R+E
74m9ExQkvHl46MhV6F2CcB2HTaT8zT2QOFHRHJ6l6bD1TfBlVdMvKH2VVeT5L2Ny
810V/08BpGjhdrl2dAovmlrGAXKlQlcyI4+l2sshUxAB3+MLOKU/M4ZGyN16jDZ8
JdhmJp7kR02XL8gIsL7Ugkfzt/6iwdQo0ktEPA0l6gL0V4sKTfjyb6qu3srqBL3i
GOO/s1xJqFX+CvOVuw1+rJeuThIWkszvyCFdCoYzMoEVlf7k+to7nYOzL9vyKun2
stSG1gjd8xWva3JsxQiDRnvjAVrZqYD96HVRqr3v5FQRPgc5qL9bN6eGsHm3y/GO
g97cBhNSCygy37YTlHy4Eowq3Rv2cMomWQNG5wi/UKXD49XEyYgwLaUv8fHY4KPN
kw/CkWfvzFvIRrXNI8LsaO++NftxwSf0cE2NEZVjm3JlCcG8x6IB4us9fT6exuxN
idHmODrEovEYZpRGUveFMoinR0BZ7Qhtkg3snpqFflG8eiViI43TTjzAx2H8y6jb
zf9G3eWI8AMtc4TvTZoh+P4NBaQGok5EyciO+iWnE4J+aXS5wZTZxc73GomHJzNi
OfOh97iCt/UQd00YTRmSp/wjB9mjpF2rWLbMnAjvANxaeyxzqftzItCBGgK18szM
KQvBLK1jpZzg59qanNuehiULDidU0AynXor/7vb1r92hOEY6VJTfBK7PZOb1eMZp
/bP3zxNuMmd1fYzLqr1Zl8oYKKV4K09vx6acI4viCFIp3E3KwtdBMk4h8ULho6bj
HGtOA6CZKFnu4Qj96bCzdfPHggCJ138NhwIBJFC7XNUP0jyYgxqgMlPGUrUeuXwC
4qiC6McLJyrs52ppbcnQsLTIu6jlWm1poEdsTqlvl8+gz5z+EQWTK5Gg7u3YTp4F
uDPDjRiagRLUDuebrdqHvORhiwjog1kpDDvYBYhI6v8qVmbB/vEnjsmU3rSDpdPb
nuKTb/ORfOTRuyg3LnqoL9T/AZGOgheQX+Bo5AyhEcz7KVMJKWApKsUdNHvq2bJG
yVXSppCSe5ffI90P/w4rk1aWO88iAkODpnBRaGaGjnB4cl65Z7Qj42Nxzh7LyI3f
aAuhQkzGcYMo5uPCwTrLulp5UqQZK+U98lOlSSpz2JQUlfgNTcSuEEc/MULw6npI
3XUt89V6WP+YobIwA3J+d9KjQ4RfWKWWE4C3hzbysfPX0SWX+z3guicO0QxTfoSZ
G/8mI+h2R0plcF0XTAvTtvfzHzQYdkiMxOS5j4fh+g6KGMFjQchEtyByDq8h1Ys+
mP+FCps/AkNnHPN+KxrGbGi3XFtnqJJSBVwF/l3BRqlIsWXYfN45SNZYk1tTkxcB
p2cBsnGFKESg7J2m1VGdkYcCk3H9c8Dyqd9lQUjjW9nebDK7R6KUFX2XCPcjTLgO
rOONbQnDkn9r9jMJDB5rANfx+1Iorfz7VPOaborJw9803KpuTwkV+G6WI7IpCOdz
cqunc80NR9dGFemd06PiSars0RG5/aPaWkE9IIPzfquwMi1nbMv4IiVIWogLPGU1
ycMzeMwNr8EU1RHYvWsSO9mzzsyfAlKOegETgLhSxfnJtb1DPhW9w8NoeV5KFeEO
RBNqbFgwnga+SOCEerdX2ZNpWI4PYdA31bpga0AnSTbByn93n0kjzXfU8OUxF7fX
yrraMc6xm49zzS2vZHwGOCJPJ0rQ5LE1ChedpHZpTRb2IxTUgoiRIKGpXnc0VR7e
TfzFATYjKCJJAHt6fZF+UL/R/H7szQQEglEfqQrLtIT80G/aFShHLGCFAWSUH60C
OWd73WuylKXo3TRcqZL57VHZ6TPHchu9zxrafBYKKVHOeGpcml6H7sRIIyql06SB
Ao02j/rjmwXVg9WbQo7oSmV1imYEEJaFO3FzvCbPYyrzPsIDF+jH95FYLa5nktFy
dRwYg6sGEizR75foJlNLhZPvifhn4K8kz8Urnq4fLZTyzObsG3FpEY1Q2cbdbBri
29nGBoeJxnuiEg2LHgEe6aPhQMrdXAXwH9QE/myXSctYoKj7IrG8aIC7jDyWnDvF
kjp0Jj6kmwapTbadPRDgp4sQXirKqf/ujNE9KNqfGrLgsI0iZqlqwezs4hAESMzz
E8Ja/wCNBW5Qu6LAiq6HJ/9szM8e6e+gMmO4YtHXP/D/UfPZkMbZB1FiL89JTDlQ
/Zn2bQD/BC9ZLOw5ijTrzCgJnu8Zcet+1tr2nOmwQ92Xb++9Za/66D4ICjvl7Cv+
M1hmPY8ZeNWv0OBa1tJcAiXGH5AKK4sS+glRbT2wZqgPZEsxBplDol+YWGF08J/q
kdmA+GsjME27L7Rbt6l72mL986S5Mq17GtRHCRgd//MCTAAhBQF0PgiZXIdVvdB0
DQQ3mWuepKEeSDV3SVqzfA1+ajYX+qUJcr7S4cGB8FKV0vesMWGIpAieS36tilus
bRz04XcPhLR7LZvWQZr1o9AOJ7jqaPOeuoLkbpQEkvLQR9eIgwM13g+cppHo7bG4
6FjRrIEncS15C3nn6DUn9iI55u8DKNSp1h5Sv+LiH9g8Iq9SgwMtFnr1XiRJ308U
NQMe2G+g/MfXqJyL3yktSKzxs+3wLr6AkUvo+7Z1OA8hDvFetNWcnqju2KKokPGh
2y0pWDhYjhMY8m+2Pw7kzQLcGihlbNVF/uS7GWmuMBFmxlC/2qOL0IsEFQ8IJ5dg
epDIgeyFGvWFrIbhtC+ldZinOFqoCBcv8z7V9FL/jykT0ihMadunaIPGscXxhz7i
ZtEw9gh2XBvAjQgGZ3bRnErhQ/4LKZuwkbZV6GT6elRtZ0vGLQ1QLZGCnmW/gEPX
sply4PhBURKkbEHVWcqgiweBP0UrFOqgdqgMdpeGHyyU3Yok3iEmGBzIzh+N3ngG
ad71VcV2kyRlRiN6ic8pq22a62YGRDbd0IBjPWDJvBYE5aBKjk8HBTTJXVUbSqCk
ShsGFTcvao4sZpN1BPWOC/uYbwOzY+1b9R7cjkMjhHjwalYy+DtWhXONyF8VSDwv
gQN4k1UQkp5jZagWJ/2qcnJajYnRDWpFzB8GEpg0owb5X8+4TsMu4S9n04zvDVyz
ocs4w6FIiaSwlm3QB4nwmJP5AzbvpQ1WOsoZSb4g7LiG7hburHjZf7IQzNk56g3h
CXTHL7q4WDU1coPcQ+ukMMCLANUZDZHDQKI9qAxNljEUyntqs367T6eg8mAF5H01
MNtQl9xoouTkJbohYMTA/VpQXza1pI3Uk2zLi7Lbk2Zw+ELUomGmnUZKn6ygnsTb
VNttQYOUpBvya22qrxiC5DhjgF/w81IX/hVJgfNfusahurvc+OAust2RxcBWmhdk
/XDRp1vDazWfXwn734hUh0+0+aE5bPyFKkASjrmLqrxOB87y9bKSyqJ5uacNkCz8
MrMyh8BwLnYmgVkPjjezItnzvlKAsc0XUjVvwdefnHTP8l74bTnG4ztYb2HhbZFD
FXTTHzAbpAtt5la+FVL96VB1OlEPvIxqZRsaFyF2bKdmd+JGT6TrtShWyv1axVYo
HUFbuyqfn94wUL+J4JVWeAvZ5NtHr0VdT/VZQT2emYir9BuDw8JhJ8noL7YLGWf9
SkSqos9uCRkuKNb1WoXo7/Zu2ZKAz2PriW11SfDlKjedZt4A1qMyA4FD9BSPZqXE
0DcEcmWXVExucLLduKGOy36mkPo0kNem6itqfiQNrT33FPaMo60tiy70rTk0yGHd
/fYmVfZ26/uU6kOnY3uYXr0QOW4HzHcTgj0KWKCG49+BgdluxdGtyHB9zXj9KaXJ
f5FC/LFCJX+9QWXg+4rx5754dLnNWliuviCoigs3bJ9Hjt3Fu5upum0riq8VUkn1
i8UwtFofVEK7Bfafw0DSYetEYdM17SJBdJsW1xhN59o0r/yr4S+1g/06AVjEwxdB
LZ0/FvpC0/XiLQSQPXTuyVgolMBkxU2ScV1zVtsEl74KVseCLhKsWbwWBe1OsW7X
XtP4e6x9uLRxkQ2f4ppt9reAtKTiWH2HMDjhD9nzhsVuHuT5fuuIJLrr22xb75lf
n80rjGM+KdZQplOmtwpSkmWvEYozzXk9QTBKiVv/9xrSpQ3JqSfvKySwMksEhV8g
b0esDbTDj3A/UQ+P/MsFxo0sW04ByYV4YdjZIqecpk9HonvwnsY8D0M9FN7Q14S8
Da/qpHlz1oH0BHoafa0B+XtpNp6T+I6YcnJcgayT48VFtBcfpl7rwHxwNoqyJGTX
FP9tMy4HIQNASXNopHu1wd5D1lIh38nInFkjMjHMnOnXD7Bszio09v7+tSOJ9opr
Fb5bHhVz+XGuk87sYvfU2rX2GBz+gAJXl/T1fvQVDAFV6oMOCNWM+NliJTMqv0nN
BBlklaKjUmWYHXD485QUVT8/U5xUiSFNGw0zd6uBZFUiY6DM1DN4DZNgNnj28AVM
JJ2WiwBMEX2HJCdai//X5sJs2DR0lxMMV6H4bGlO4gpxlu7PoGiZIMlqNcLem2q4
9vQftGTvt0j8aVNZAzKE7qDC08N0paletJry3vlhVZTJ7ACXB/9XpGpDqj/xvjjG
Ti3rRiewtVroJcBhcNEe8pXMGHY3kLy0hQJIaInAEyzD15uV34P86+s7Gf9rkx+c
7isdvKMeIWUBwCRpGkozi3TpdIta6TrBNLdQ+Ypd5a/+oS0P9GfqbMRPDdfpIvKt
GxwMKknSR8cYvzZwxrneUQpqwekBCrEFTRsRcdAvcT1ig97Z3lypCFYDnekSzRR9
su2yfkdZnxeAWdyYA/h9TrVeSMLXsj3KSBElkJUQxz7NLNXjl1Mq3ukPedQ+z4yy
si3NFOaUKxcbydPys2MhCp/HfLs4Mziugq5fRtyYV3WS/Budn0sIGG2EahH08MDy
OKqDVDZiP6rkiVqGY441Hnh5ufm3zgJvySTCcmKLAYN5x1cjVoVuFLj5NLIAgr/A
Z9UHjc6F778YwvVMCDn4xGdv7IYA+NQQWbhyEJ5GFJD3Q2cYklsbDRuPk64iRp+C
sI/hl9hzhiIl/Kch6ax+y5wEsLROT74nu78z1aTRCO7YvF7A4aZAINgh9JGqtV5b
xvNWemRiRFsUR+8A5MfvNbW7N4OGNQ9OGlbkl96o2ISeYhNdN0Y1FTVZJEppOwwq
oii/mIa8qdRKfeerP0Y89tvORzzjRcCMw3gc5e4rMdyZSjscLyPLTs8whXmh0h/g
dqoPhAkXFhQHb93p1y4xGSO67k4K/ea6epK9FZ7zHVlIHIUSN+Mv0j9souTZuSB4
aDFP1kHNTuf+OGqfRzOU9JTUp7yvNIp6Uv98mV5wbHimDuhGea1Uyc5ubESfGm6l
cSSTnZhoRZ8cnkG7P9RgFBe+ATyuSnrNHbzEZCVExWn51EU2ZMKD87dxPXLEK3LK
wXMKedCJU3Z+vk7ra2SG/w80sy2/DTsbGqhpPhTBXHwC0S76VZsiwmFd+r40mwUX
8v3v31+V9ABqSNSck/OMGKMT9b7nxSnTmQSNpQtLGNmzocVb54jSsiEedINI9iRQ
Hva9StG2Xnp1bHbna+7BLM0KMB8OfjaQE1yrLbpHXsjeEaUFsmzRwbegFeUQ53lr
+sE4VuGGjJSov4B9Pkl007tVmRqGxkXOKK09mTmxmrvP159hbZDyL0t7bPGangzU
m5BsPOyNT2JcqOInAwlYdbtxCokt1+q/xCkEXZAmj4DDZw++2SD9ph7Ta4AzBOGF
20jcjXnR+mrYTQGQ47DRUAbvNh308kuRgt55en42iB7onkyt7Nmc3CHMx/hmziEe
q58mXnJ4Aj66UHbheuB/VTqddkBOfPR2T4h3HteMZ5CnZlX7N6i3r7yzwUu57qP9
EIywqk9l8HrVC3n5koqs8DIGhZNOsl28s/a3sgM/OqvXpZMd0kjYJrEavV7oHvof
obJ7Vk1Ee+iPnuLp6Zj1ZGsltXTCXdN5xQ6IHVj+6g+9ermoLtLcsZ9/m3S6CR35
uvlbabFdQOrHybSIbXiro+gjMNh/RMTGS1ToRxb7Uj9755j++jtlBXZZFLP7QiWx
sEhhV0Ye51+9FUdfiGkcGBuiPUybWXvRmhQFcKezhmq0xrAYt9YR2KidPNqX6L8X
hTe5tr+3BJDvdDpE8TkNTk2etEMKS6Gyr0h39VZ4wYXABYDXUoQaplf12PW6zxk9
e04IOMv1IyQKwAqy5u76ILWX77EO4qkO95nnrmmss68LmATQY3h5y5rWRaW+u3ly
0lPUGYFtDQPoDR0F58HZrKnE2Po/gIdD13LD8guJngoCvVnxKTf3YMf9IZ8ZacES
4e++ROBzkjVaIqucQqe4VzAqrbMkiDWo8UaTFYADZMWgxKXzDuzkQCaVg9d2dBgq
TIJjs3U4WneF/Fy9RluI0Ve1DqPDAyXPUKJBQTH732Cx0nzxzuqbfOkqvZinzKTQ
UqHliYcJZHxpMMAnJCtPNe4r4ejzLgm0emkfLB0mZOUJRFLk6Ie/QrbeMS3CpT1S
mGP1VeGijWsQ+nX4ILEjConJKpP1WQVrJUWboKvcetmUTt9lxIvZO5fLFA3bVW/X
PjLUdvP1E5iI++ln2OV1a09ZzUAdcufyE32smbZKbGamysh8Cn5CfhF8WhA+Lk/s
l6CxQhF/RuWgzfJ5ymhCkh8TxTjsw25SR4DvgdJtC4adZ8GKuKUR8P7oJJjPeHo+
Dz29daSJFllLRG2rZJrJVowsXpHY1iE/hj2oR6iuNCGFr+MtcAcuOm62Uer2Me3k
AQrF0b+Ke7Jc2UXXnD2BKdtBxUQWzYTJoowr9H2mAeUsz1WbJrYNsbyFH7+nvwth
0QmKQy9xu9fr9sRpnbJTL0ySRedyHAla25inR9ou9NM31nJsWEIXASmu/NeKosY7
VqsVuatVEOF/Elc8uL3z105RJtO/Vuj5ck7jYxr763ZKVzgigFbPmuAge9L4PJzr
tbPeT4toNYw4PF5YZ+0Ti1Pv3W2UMWeKWVrJr46rXqL+wkA+i/eIYJ+R6NM0balS
QzT3RBgkmO1UFXsm/1sechE3e+JwJ86vQnL6RMgZvSWRAX1E7XI98kkFiMX3LmNO
V49ZizF6QC9ZUkCXAkAu49vtFk+BZ5d2OtVLxobihopnrFJZtlgzwNgXHXVWH2cB
CtUMe2/SgznbxxH6cJUwEUzpFip9MLA6xprnBaT6DiavhGiNKnpaK8hacPkPQ1k3
EEULHy/jANdatLllXmF4xMdt7eEIPRRH3W5vPIsVv04VYGRzeSZUCsijJMQm6lKj
cZ1uR+M/nTuUdOz+MQVXa8BKdAdjCr10qagPzXm8s+Os0CmD+Gq8ARajdXUnGWDa
ZH/T69A0TVWzRFfkNjVgsngyo1En6+n8BvtX9O8BmvmfciCevYMd/6tSJsyKYxSm
4d6X0SFYx42XEq2ggfURQKFxEi32eirviudNY0rQYdd31QcrUlJj2lndDCVosrCK
qAOWYRaLVSEH23OWLPftwZiFeETzKR+tin6Hhf+txQnbAkYXAkB1LgN7Cq5AQ4Kg
Xv6idldTq/NXf5uQFKzHgptdVmm0NAM4bCnPl0YTs3ZdV0aWcjbOIfhL+f/VzR2H
73GlUIrEHvE2rBTjyjektbp+xJHrwpEK1RGYzGdn8wx3FwHHp70NYTKaHiVuz8l1
zCfFTAzoOiWHOl0elcCOWzHnb9X2LwC5IlM1wbYjd+TFMwL5Y64TA0EtivRKVJCa
fU9pv9BcKUe9EINn2W9En/AE082DnllryhQ96B3XmBGVtQ1C5Vdm4OoudJGnoO/e
Kzi18dMswLGONyF8nPsSVPcLaEjupAF0CzyegsQoWJ+IHx/IWOTZLfx4podOL98D
AyRjVYit8l/0/O0j/3oPv3TCftkyFWAis6/IExWw+15cizPdb5/RAse3Z9QZ5qw/
gLtA+UmpB/xlaNtUC2FgjSu4LhaOWIehx121SkuFn+yNtzdy9M/S2heyYjam2uLM
EwPZR2B3WdfqWec+TX6wwVwO30uNJ3zkwYa1vnEnJHKkRN6dGEFNf86xszLhgNCY
2yuJgQmVnBLyfoL/f7LGm/L0RZPX2NY1cBbl8fgTHFdK9jIdXgD5Ra1xAOEkDo08
fevtm+yhjgHR50BSHUZpWQqRkbIH87fftjM7xSIb/kr7THO1/bKsWpRU7o65bEdh
j3t4j9RfOS++2D43EDbI1SA8ikTOuUNiTU/B1Dj3C/T1q52L7OxCdXd2evBfoFTo
uL3uYp78L3vXJNUW/W0Avvd75gBqz3qLOUn46eSyQycfcYR9vAL9vHR9U3y2D9nY
7GHVpaXLReINRRlQS1tFoSiCFJYfS07N8RnFiF95Gn4b84hZPhwwpPG/oBZgQ8VL
siZqcR2rt4LfjEXmyztt8mDjosdRuQKrYv8ND4oR+n24TyaKBFbRvsxuU4fLcs36
L3X3yuXcAK3wewQKGjaw43h35+t0DEeq0JEq/gdbN1gYnki8Ie+E753pAtdi3HmT
2C5to4Ulcp1TjzCzQeBBXWm48siXaItGsJYs1EyE4AJP+ns8hfaJmNmzqzs7ddEm
zxUS/bqoZ/vFCZt7L0OPHfLDywCALFdGhkiEXlxeWjcM8enmZTp8RyFx+zWRmJ4O
tWxxaQCqLgwKlGeGo7wOUCv5W0YxDeFe+guig9CCt5WhvjXZjbc7WVwqxpLupQmq
IaFEYt0BNzlVMOirBzEHwgpYSB9fqXBrFadY3NBPIM1JerdMAaVxZRD5eWRnU9u8
2e+YWpvfGa25NJYyrM8m8V3ms+FEnpf5g50ADRfPM5PodEgpyyasd5AT9JsJHqAq
MM04N++IuE9GhOX3IZkVt8BW48m8AKcDoh+3sfUf32h1HmQaKjFD5P2/ymD7IEwW
0Ajeqr6LI6G336CmvtSlYXRaJ+4Jd8uxG+3LI/w/bbPszAPpqYEluz++BZq+X63u
dPJe0OFHn2Fv7CQMUnUbmSKSf0PMdog/AH/7jj4+7ddHm0wQs71PbazVqutW3NSK
i4CBA4j15NBYI6NykeXXYaUjvuGcsc+6qrkE8kkcC5O+wpMb0D88xY6FtiEOny8b
lLyEA0cdkPf+38u9+/u/URIs7gwWogonduAtTBzMZ9s00n4XtNenS/I0IN1XYvq5
n756UlFpxlsqHAA04f6pzdgY8fGoJ673rZMN/o4AGkou8eVhuQsyGRKwb8WpLLFW
uTq19DAf9l2Cg4Q+TXtpF9cu8oD3Op8Pu+gpKOJHdwxrVrpzZA8G1+mohOKh3kyY
rrqeupIx9kdmV/6bpgQ4x8B2548VMtF6+8W0OMpYp6/YbMHNlxitp+4RsYA2Ve1J
yANiDcHjWYiHMHy2Q/YRJshTfePPMmrvdzBgLENJyfpGZRXWknxLmKf+s4JbB2xM
S/OT6ugDOfurqBPR6PI+lVq6797Pz7DdR0B3wDaiuWfgXLTcIybs+uYrXqN1gPlU
FkXQx8Pza2JG6d66B14j4nnAvS+3XJ+jj1hRUT1mImf6ja08niSjzSqSEL8L9Uks
cJF5wySnz+b06FCZo1tyKcSAQYQ+fS4GNvhgY/LxthtTK27k6r+B5EpV0AKYSt7M
Zj5zgjiooCzxzWzdoXn5bidvUIzDWShGuC0AiESa4yB0pQXHh4GZf3xw6b2GP5Zk
a19cJHdGK8BRCzUimL0NdowoQjVU6jOFaEn2twtgOd3+7gSYrip4pLIQc9YjcBBq
9+6C3qmbPYoKeykHnHuaz6ZD16aSmXZE9cTNKzzGaXHarg2lTW/TTsBRRX7Mgt6z
FFWUBbMaf03bGniovofeQ1KtVgrvns67/UUmwO6RoO3qtzfFwlhKB5/pMX5iQugY
NC6EeSZnW+kjrRu72MNCA40TVJc38gpP+y3i+1A/LChjLxln5bFmG1JQEPOGQ6eU
FBB2Llu8IJ40T24QPOeVw2Sus2I6bhdW9Et//cNDOE1KaS035fUDSINNgDekwSwC
YtFp8cqv4dZO3f3/H68Z5aJh/kevaTsk/do5O+Y51UpbzEnlnnsHNI+hfMk++VWU
lECyL0vpsX2MoFZV86i2WxD2nnsiYz9DeKDXeRh71LcwlJVQlB/nqR43Rwvoeb2L
4XYnb4M5cCxFCVJ/KEZQtqiJvHWaHpemn8jpBlNiWP1BGcDYpmr1lquidQyM0BHf
TQ9GRMslubhhkQBJ+y6bSEoQNa9mJDHXcT4IPNndWMWWCmXzU2A4mxdx0O6XL3vX
mM3BvxVAYNG7Z/o5kP+hVubO9vosi9sFUhcXLfFgsEafM+E7fGugZyP/TFaJiojT
pmxvfS+E3FzDrMD/8EHYnxOdn3B7zSEmScONwOfwTdQbzxTVEqZoD0/noHsel0G4
Hq+5XsPwGbTfKT3ojMIUyh0XRhKlmmPsqiyQkwj0i01Zoobaqi5JXYWw/hWVqObI
fRd6E9orO4s3+BvXK8RPSrVvCI8yOIzSmfpzUsQBEPj5E4Qw28wJRPEXqIV+1NOH
iF4TDjFNlrUGxWlI0VF2pBQrzv7XIlXPzGuhrHCi+4sssZTNJcWnTk7cNCBVVpWt
ssKwB7oDzQZ0Q7ZdFE9Cyu37MACAuJkQL0Nks9bMF3jOXzj+ZcKkQtOyIUszWIfs
XF3Njemtgqq7AsyMOulKay7b7WZZZOOt2uhYiMHz1kPYOJghbYBquW3+1mHluUZk
cZ0t5y1dGrktuufuqmDWfu14vtdQ5Sti6mkeeSIPbuGRBXHTp3hApdIX8lZmtS+E
ZZsisL6YIo2ZFQzfEcwtplBE1GjEXPl7/cuww3w3aL976pZIKK+Czd2hEBn/r8M3
vofSZ35pbyZewgBwUzzRHhI5tNtMA96sJKXZsuomO5P+6mkBPP9WRAlylV9Td3mL
9egnYmMBtLBz8I5HXLXX7GToA06mUw/xLXekz7bVK+la4XRYffRHY1XPtlOc82eK
etFof+byyVVAaHi6D/5mLVqZzjw+3YhZM/qnzFL0JEJZI335AnXyOLI7YHRZhMKs
66xQ38J9tHzT1udPAEIyeAwBVn+3ssMErmSRX+yOpJJ1YzoG7+nDp3FFZdoLlF+M
zVNnkcMuP4IUlDcjQFCO0MAWdUYVOdUo9DG5IZdwWFf91iEjO4FwT0jvp6oxfwDH
ri8jjALFl5dXs0bT8FUVmvKAOdeCMunDYN+Pp9UjkGnrQDr4LR9Phfu54LMagMXi
Ax+irXI5Nzlryl4OE+QkyZNw54Wib5PXMbPFCd7N4g22UYhYTvgmUt+pqH26bwXs
6ZShBiEfPaFowxP0urctzED7IB7FwwzcM5lTIxHD16hVRMq5adzGrdCwNTX4PZIy
WqBuB6TsGbdZLs0E0R7kw9Fsy7LU79eJS9vGDn9XmeCg6ln3ZfwY/STh0nvvF2F+
qWM9myL/jgTLUbyCiG36Oj5Miw2OlM0veYWc6HUz5554zzxnFrFsbaqVeQFom/di
KZQsVD/B6bcBTLJwm/Z/9u29AwvGMBCY1nHv3KHq1mPhP/Zhm6DQpmpmJzgq3Egp
v/tTzSKMVcwobe0AAF/BiHemlTTfSd+zzsqk7uFm30YQhDLlu8hs6S0fQ/hyxEAT
1HyCpHMecwNodSdaxgpf94K5FqrOBC0Ks4SN2pSqzl+U22DF0R21RpcQRRg6LUMI
CCIF/xwVi5uk4iPmHNKGvt6aMKsmyBECYiKR7mPbJrrH47RhXYlK6ciBtG9zzER/
Af4V2RN/eJKbyxsaR9Zy56S6uONP8N+VMm2WeQifDGYltaEUv6PFhRNrUP22/lGP
Z38utR19dLcDa716rIjTy67QocnngQcUBPCaTPjQ0D15OLBuqDm8QRHDIprixRBt
+MVOkvbQBYlELJdlrDAwF5aW83+zSJeiaEsTREIdzqrDrRmUaae1n01npYpja7l/
xJqIvi8SJQ/7Bh2EGr8JoIgcl2RO2YtmDwvtotKCWvjwxdNYtvNJszrBwOYr73y3
o9+RDVMHKwm8zWWQvFb4Bg0m61wNgm8MuoEJrlcoQJI3vNqjc9C7aD130P6xEiMj
/UKlo+12xOpP0gf01zdPIqYEJtrlcpPaVFFfzFAWlMLsV456ZVuvhh+9MStMXuQo
NjqXx3oCmeYBAy5WnVrRtjEZ5+oD+dseex4q6bpzJisSl1GKhSO0nt7Np4qgAQGj
FbBZwcgWy8Up3gaWfI+JLpkYnQU6m1iYxljVvUFFsVtGuPfEAgWVr+B3EY/rX2V4
sW/oZBlSamNdo84fS+EGQk59WfPZnPFd5QZ4cIVAyH3v6cA/+ogPDZe3QD+gPOax
JyBfLsN3Gw166jrslkjSaLERM+SRl1U7ZEuRQi64y5OGkmksO19KRFoNulALBsGa
cmmESsBydm45lT/On9CB/HdM/C2ZvbaTYVN7K9vQ/W+HOrwskgXZhHLV4T6rmOGp
16k3sRszIHqgmHHbwidGIHPxo5YiNEcbFWbNY7wB88/PTpVhCeWtnejOf2nbwYk+
TfzSABIPJ8yvZAiRv7MSgf2+D/zYwMPnp1np+WbNsYttoF5x4cGTsJ2QKqskRp4c
X9P39vH+Ubs5pswiGe6352A2c9ma6O1XnSoy7wW2pWoCEMIyyYBhPlo10QNBR5+l
A9HxwC2bVWy/jOWmJxNu+EmPy1nQ6+P7En9Mc5l0+9gC43DL5W/8GRkKIZId3P76
gzebZnbkQALT8448scWU5bz1MYg95GcdboFiSqwRIHPOtZ//q9u5j73bjdZQZWJE
XNyMaCvZ1bMAQHmpsfP9kkf+Tt7xhKrXtykKzD4wvVBA5wezY9qwSMaxw/yIl9uO
F530CHh26gg4mrcX9taePYqfYAv0qq8GhN2pNKiCI7yuUQ4wX7JL02N5MM2QbKzN
u9SjJy2SfNOthUIxY/wGp2hTqFUl27gGEOa0VC4oTm3q/uOxDi6/MFIW88KBCx7K
f1DTKJmLk4Gki9jhcPSnJ+J1tQ6ARGWUsZquk7vwaRHR7xXZsduqqFyXgK9LTuZk
yTy8+lUif4E9bcu3sDUjfSToei3eG35ZtEq0VlfJP8Fxs7UujyJBI1eOmr5cUok8
4bkuw9jNARRKBSe2Qwe5yPwOcfs5GEWRrohj272TIndgdVYwcW+CVYvRmuttoEQr
U3qx7vaF5XQJ+xJ7nJQRRcmF8dzXrnJNVSOMEisGH70uNL+Bzm4XMVapcmOzP2i6
jYMtmHa45xtYERrUydqKy0r8s//L1o+4xhEDVQmKnd8PDNnlUY2xBFRoaEdlaf0/
KTrCbW/srjwIg/aaiZbcaCbDPR9e8SIYRWDEzE77EarAFihAhVoMTj57UqTVnPIP
QPY1nU1JPfVm6vGpkj9fiyCBNjQQpj51HZTLhkO80MKeJ6x9WbQo5tKWdVTv7P6V
0rIeh0KIXDrX7fHGYEV4N6g5VEdGDR3/vtCqLDUj1wwHHA0IbLmLzeYzlZ5Wq8HF
uwkSDWFLdI77qgCaI2yui44GgqsNy/4t5YDaKjuoA96vbDAMFmwFSufKR07OpFxE
DgKQjNKGKQYRht755DUKXIw06sZRASpoEeDjwZCEoVzx/j0b+3aNS+1lDSuPmClx
/0spd3JHdTvloqrRuEkAFxa2QD2bcxWtQp7mv5b6qNcF4aGmyQNiLr9hAm7YBnx/
/FbQsTFaht/Cg3QdXv0wV8eO+YvL6q+wqxqTOfdLRIkZAjdpJ7/95xMTrDr6NPo2
Byk4zj60EpC17MyTk2yWL0Or8ZkNzHr1yN5I535xAnokfkIyfych/Sg/KCS2JNI+
BIvdknagzVIMeMj6diU64IyKZqFJXPdeAviHlAOrkv/u85IBchBzNafb7DaAQViA
CLiFlpbGZB6XNP3sPHCZjzXmqPka15Phyo7HxUU/dmc46gql3k7agpQEr5iAtZa2
nkslS5X4yLrj0bgImuPoYbs1MoWqmB+7evTHy4h5QFl7lqGqd2ZQX1EUe7uNvVkl
kq3hH4J1lMEG0DVkB6ba2FTcr19Vr8Jgs+r5nvdOWw3cCnmKmVmmRASKElpk9wJN
SjC9AYObZ8ommb+rbz/ZiIG9xoc3CPsUa01FJR3S3vsZ2Ij/XKD3IXXCjf6jbrZG
VLlRuZGz8dioiVoJdGIb1iWPAM7ZjunAfi0qa41RURaWiVXqV5L1Ik1bNvSvg31F
NM2TXMibOYHYwKPHI93ArSm1qW9F9oze/DhfSRarZU+QZzKSeWELgJR5jRLhC/zq
dNuAtDE+I6hgUjigk3Wr6RMzRUB8pHs1QrvepHM8X7Y0jK7kJfVvDXEqrQT8FkMN
ZvnWGTDm/x4oUnENMYz+MzrNP6UzBdM+M9uJcNcmmE0w2fZG6SnIR32+Y5a1eHcn
DQf9iUfpK5gj9Mxn8h7QiYwvUL9LWCgtHtXzrrN0bKQrU6zU25JKcoArVT8xrnlE
QZOuJw1pASgVML2/QVk6/JQTnHQ3zn4CJHWskger4fB+HOPIUIxr22V4S2lRdjaj
o+KCAeZxT/tjMAv8AOU8+gKyC5jmfWgyJacWRdghCyRACZrK7k1WdDKOCqoczWaB
poZqZijc/Q2wb2KPkPM7b8lyOPm70iIK5Y+pFBkJL2STlSljEWEKrByz3tr7fqH4
37lUM/6A2+hwOSVxLbmGsN/GwL4cPL3gRXToHKYtwCxNFMZnUkueZS/Gjkcobm4M
NJTzTlUBoJYcyTDCzTfwY9CFbj/cP5sCBUIJQ4B+fGJ+rEv5Eeky16+tmx0QYj3M
LrfpHXWEZ8R7CbMlUGJXa9w9nt702wuFsA6WBKB9vsJILwcKxwqqPjTozBUvPtWf
G9+BEtI6b3WLncVDTMMSATbVbFIjvyw1lwnVBR5CqLFDzNYH/Ujo6ireP9n1rMB+
cB3WyUOU+w4hP684mQt7FyTlFY8R+cO/q9rtqk0XQ7JW9ArQwm+bwmhlUYySXktK
Dl3yOcRFnm7m/ejRmZD1kHI0Us1Fq7ijzygk7+XCOGFNDi9BkR1oRv0/WTFypgdS
gxXrLRv1jdJ06JRlD1mfDQJSxH4IUVR1zq3JGkWXzEQZc44vdjIQigO0ApshfpWK
sTpWGi6iiaMYI5bSgQynB+B3TT/owoHpsGFxMSk3v5/AW9qBvdMMZnUonYgvJwGo
I5CXhtyQrGeSHtZ4Qe6rFpINtcgvgV09pWvCR/coxCoIVXsuW/O2+bj8k/agUqHi
WO1T4fYYBoA+84HhqEJhYEG9coCGNA6ZxbMdhgB9TdRRzREHWkFz18tNCq9xbWk+
HdBgQrIe+M8QuN0goiTQMrFuanJjv0WN7Qfg7Ux0NZXJnKZT3GaVWQ1ERHynPHki
bGJK1VfgF/fGJGmLqy+e663CIPogF8apEHPo6otfH7i6M+meKMt6xAi+pzRyU8Bp
Ma0CwQeFBqVVpMMgle4am2bvfCbV1n1zbBDRrTD1cb/InOmxaNptD3Y5O8PZIpnY
ODSRUSg5iJqktRkzCGEngnTsm9Xht1/NMMj+Hc6i0aKzvt5Rmzj8il14gI7zFf8Y
gQ6lBHTsWJMrNQTLXxWovYgY5mD7XY9fSixDoIj9rj9NjNKqRvgCzPAaO8Ok1XHv
O7rPFgTgTKZMe4bHxTDeIBmI8SGNv8YgC/YV/rs4i865QzEQy1c+8VEdoZ2hq7HF
1WxVQI6vfN3FMQxRuRKLQxj+DsSlO1YVpXt6WNEzixUvj6ix9Y6IxEeNwmnJWFQU
GEMFohgeqU9DL6hNi9UBMh4A3QB3PuJnWUwyls8d+MTSXIWnCMVFyjdMBhT28XJK
jUJvkYIULXgDBilv37McyagFoBgCbMkBqyNaTvBLtvzHhVg2Ft74KtZK/QSP9rAi
/JCS/Wla5R+F1IsLtyi3Z1iSYjU2LdkBjvmZHDdh+veTflPw+h4Wx3skydjcXx5g
9rmBSk5+pOY8N17BbswIK+YlRYkLELeoa08InvoTuZBnPOnVeaFzz13GR2lugLCP
04XGDG6CXhRV6a7chYBdox7pl8uzFOs7ICja4vB42ALjGXFzVdUlqtWPWWzYMRYO
/Xg5Z1mAohUuHYo8pzMPbz3IfUiPXfjQhdEXVcSp4q/X1gqw0dG2tWhXKDmzaujj
kR4qGsr+1PNyWblkfPsMevjaWUN+gNjeY6yw/oLhWEzJxRwdIQAkc61aG7Gep3jP
yVOEEM4aZ4aWh2Q03/j2o6C2Kw6mibocJBPAf3WkMsnPFKtHUjeIhrtRgyKr5qSl
1Gnl10vdEyYTawInJcZX46U+Ir1az4r17ynYKsG3D/LTseLSKGCZjLoP11gJR3IQ
P68B20NoDQHCnZL1i1Jf6Ls7Gj4CVhnK3WCrDhsPi07XNTvUiyY6P1O858W46G87
rymxw0/M+qD8OYmg0nKcJO+ZXfRjLDlLsV+DVmfmbr0llOhJcie/glRRFaQpslJi
Cl4g5GSxbb8tPB+jD7F4pU1DdHcfnzWAjUebh9UvyzXOQ+NcMZpUAThAR7xCgx1M
/1q/ol+kcQieO5YHfFl4Mm1iJ+gRw9r5mNfBKtdQ9NnHaH1zqEReNB5tjF8mofrD
J6JipxjFrNg9qA/U4CBdfrTeGLzMlNLMCZHLSo/glHUhDYI9FSMgUUciCultU5cd
NkxdxTAK8YnM4goAlDt8UjVUoHEa89D3jH/Jlj+zsm5vnGui53WP3eW0Eq65IaOJ
neRvNQKZq6Lu9DQxd9tr9Q65lEVU9o67+Z1nosEh52nb+WZzg7T/Zgl/I5Ff9oQa
8zMe80/M80TL2Xoycpm2WGumBikvccQFye78Xk/i1OVvQBVev6cHbs7zuYWhJndd
zSpyvPKKyzvDsbxeU9tpM0NaGxCAHjMj/ZvIaZ5AajHoe3sxMQ5G3loKWvpyAZcg
t3wofcfwc5IqwUlWYMPmq9/7XWEJHkgt8S9bOjuKm1nvBOdDOkdsSiI5Lps/gpqu
2yeY27ycwh/c5sS8KpZ/vtbrPO/Ufp5J/cdfpHnwa6CqS8oum1Upx6UXq07N7U/P
Kj5FHPR9DCjOROWvFBCO/aTAfJvUzgXbpTENSn39orNa20npGC30pwRXvEx06wRl
SanyFP1ldMk7SilBuKnGACOPZTADjAlL0C7EtnLts/POc7MJFrDFY7iEJxf9g10r
zgJX/cnHXf89L+cL9FkKLsNjGVuDqSMJELA4vSqbVj0Bx/KnQjHPNDDtOuNDNKRS
9k1nWQgeztt119VSjYq5tr7eQeK4xbE5riB7Fu+0XrtasmZbBBxydoa3ZTA+mfij
aK11LM9im/axQngrJklzFTa6427jlg2LGvTh26WtmXLqoWc38aHBAMfoD/6SO0Wo
J8eLkcPfaTPgbFybrdGw5cJhH1H/ESnhL+3a/AsT9AVdV+Cve0HfBGpLvro8++fg
I97Y4LgrCHlbZkzoKA9Zmwun6XNCdJWgKiBZ5dz7W7tnnpaGvPw21Roy6XsSmHHV
TGQKMdH2ndbBPnXz8R0kpsKSva7isudRJ20bR5saGJMLorR2QwCsOMyXGFYVODqa
YC99lKFmQUPYsMeGn7NrZ4H/QG/fHCLqrXgjhgTIITfYPD3qEWWOZk8QHCs4WgO4
0o/xJTWFE+BfEcdpGV1mDVvlj8dsgLptv8HbbeCDuDh14egKdneLXp417k+/Ybiy
neaNOO/kv2n6YPdedtRZ2MlbLTpLn6BhEeDOlJ+3eT0D+phGRUz29EG2v6MjLwq1
Kdfzc+B3Rs7FAVPdqNY2+knI51f/Ybq+YPPJcDOLuG8EpZ8rO2K7GMcDN5ghxq8z
Pg7outjtvfwmioD9SdTdOdA01ah6jLyyn6Rh5CLdXKNWXo+HBV0w06ImJarxDWSW
PcqkhYgApxTnsAwflO1gFpzDR28LdvYlAJQRT3D38lbUWujt4bv0x9gWiXxKJTqZ
FHpjbk6ZG/oCA43OmlYEFi8Vqq6Tahc/LUywUcyzPmi/JciL3AEp5hJ6Qk1FRaCi
Ci9/JFcIqMW25ZhBlQjx3qxpZfI2Xnc8WK4LAQdFA42d2S7w7QudCezchQ71WNBP
soug+VrY4tziJhHPQIcXgR1Tji7t3ESvqalL7GyEhqzf6XuyqfCZasf9aBrVwQWc
BtWfgcyrQ683Ek2Eh4d0kluluyS6HdOXbusIbrmBtJ+yiJuEz+SeYQF9uBCdOPbu
EBJDZiTQi9Gsla6YIeDLNHszm9Bls6pqhrjD2Ay/rySdrYgpHohT3Kw6UAsXOnDK
m/HBZOMTrLKFj80lZHDA/CFTDyhdr/SUdPDBlJ4+WY8keAUkIEg7/+J3PiM5Xyf/
f3XsTQAlHX2dP4+B+Um3bAzMWgtOhrUgMIX7aPeiJI7QMTLsuzdisq7QTSSHXIRv
6BQoN2tF5Zbku7iyx9rWHAVZZyexSf02ypJzCKwvA35AVxdT4E63xpwVGQ/GmKm1
NkbxL4edSgA3l5NTjFhDi4EJhz1tfZtApQk40/ABV/dqAWnnn4LfKqRG0jbU45RG
1oHXMiiM06uDYUsBseds8jmui5p3o0KioD6uZyuS/MwaAheKJKCanPBOCdhva2oI
/mlVry3GiOOf1hG1XwgcDoCAMD8rUb7o6WrQj8e4YCirpJrXSOkfb4hDr5+nqZ5k
lqwJl79ln5Wamg9vcyH6q3TtOOk2q3QLjh+MD7kBlxiTCyitcGcio/cSfknX2SAJ
Dv9ca8lSAM6bBsVirIoSXDfuHoJ89yAi24YwJFqWvh6PT/qksBqR0r7CkAcXlMi/
Yq2YUR/8UmA9aLtGI11TH8KpsRHx46kbn9Zd3aEBbTHADZguVJNp69516CG62Bs4
aUV8/oYMxjLt3xUVdbhZ0H8tXaD8DS8nuBCI2x/rSWq2ALoK57aJGbsBdgoKORCX
Z20jhSx/Ly5I0aQ1mz1PhJ8rMP/fBLH1urqFn3x/oS0oaEG2MVIoVfmgzQzEH1eV
isJo7hXIVUSeaLik2LNZ6hExakx6yhjHTU87OvCMWqMmOwN/WJ5cZM+o2imrzNCR
vvrDSFPId/ku73dynaoivbc6nkBZ/U7RaB1+VN+0v+NZI3MY7ACHuSHi8O9LiuSN
Aly/vl1wehAwbyLYvHhqpmfJyiBf3jqimLCijnNoFMSk3RW2jqKjnuvPvUmSJc8O
WyOrCGCmX0cXOW0VgpmrUBB17QKNqICiXtFxQ1vx3JWp2WeciRPWDIMsmBi57Sna
Be+tq+m7vyuAwBqjMqQh797etLVHrhU7pELbAwe9e4HOgB0WA8guZaazl8833XFF
6bE9unfm4uKFAXrHHAS6/Y7j/K34ZyviWJH3tfN6Tr9Wncy5dqAoRTqvqaJqWENC
TdmLRqqXl01A87PFl0DakaZ9JmMhuQ9GCPag1sJJdHGAAUrRQKFFT50Rpsy+zQ+p
CG9JNCHatabwDlCfqzuWsOujiYO68D2Ofrz3+BjrPMgPwYvmItthSteJ6/3NiJgk
2XIYe81UjDPOsphTAcntagHT7O6cDXoiTRSvqeymzpl8fy8jDH6kZXqBfdHMrwBG
dX1G8N0vNn+fHfY1J9mQKDs3tdohjDKAJi5obwi9AymfwPwG2/NPYKJn9OTdmZFr
DpmLEfO1uXnAS5pao6TfejaCcWvFuufl36SUt9NUT8OvCC/iQ7C4twp1Dd5yv2yO
h1HiejbBG1wIA9brsgdX8vOtZimU2WKmal6oz8xTebz+Ky1YlqGz4VawoS1KYpCl
uTksCP7q1hg5Z5eG0T4Z976KGeuCQksdEjc+cUejLEa1qd+5123EqZUxiezWmmWS
CzKLy/4e4dsS1azppYs9WOLKsI0QfireBRU0hia2quKZ6m4+NAynvzKXcXrHS4xa
d/zwLVstoRaM3/VqYtY07RRw8BzHv/H6XgT3YbgxG4Be/2bQ1lRFB1EpPP1/ageD
sazafP9W1J1XBfyF7/7IuPi62F5J7cdtb+n+HszJY6OLEjqEDZD9xKaSl/iOtkwH
jA921sd6kqDndxoG6g7F46KTV6XDkvyG2GXaIYkU+7TqUv4AdFKddu3QrrJVyGKo
0dDJlAzZ9tCVztX0w2LlkgyyPMfk4qERCr8KduqQa2isjaOskydhwbsjfSjpDJ+0
2fJFM027/Lbgd+Lh2l3XJ6rtCDlJvHQAEgjtvK7AbRX6PDVa5kVH+VbDv4IxLCL4
hK7gNQP0MXNnkNj8biwEEy7dSW7V+ng+nYXLYjPV+4ZPS3oR5mVRXTRsPhm8yF5p
fy5iMp/rlL4uVigcOfcPVqOZfrZk9xosIGS4T3Y/kWlB4hC4y/r6BBQk9HZuyozy
Qb9NYrFI/PT6eqJGNK8SWcjlKk6iCrxeuDZdZbx7S1eWfhT1i/Z6VbOEJQVs0Cz3
i4E5YDhVtTZNICdMf3yIzutoWQA3s3BzFrShjRhyXih5vk4qy5W2vkaiWyVruM7L
WBl+jyb5bKtxAov9YbPvStPXv7EmJWci34FWc2aUqQV04Gpjqb2rfFHgx0OgAo65
MJSAK8IbpJXeoI05fvQrlK5hIGtvSV4R3X0ViRc5CoNk1uHjo4grOjBZJAG7Ifcx
oJik2hPFiHvtCgQiG1JP0d1Ux8Taq/0Fk+pTM7xW14IKzyEYao7pc3+61cUPmVnz
/0uj3U196FZE/lwHS4ESd7QBIetHYYkVqSJV3fgv2vO7EOY3H9oDgTotikK0jSju
biJjf2yoYnBHfgAFLv9LkjccpmAmqOD7teXvLzqOABXEbxgeAqXKp7u0Fl7/ZYjI
tD3LViMLxjmbe/J3Nmk09/CwGqyCetAjcnrzeRk9kYL2lwKosxL9ZqgEhC0NS33I
v4JsRogkS9GJeAkqUg3xE9dwHDkUjuKfDNQMdOtut5y6eqNmNC7W7wu2bhmF5EUj
3dEikQMfw8u3IgY3ni6vi5foAoFKKj+rwJ+YsIlCLT1lPllRHJ0CQasVLoZNIe//
83LthVufbMUDSOKewmYUIwm3hGnrO6biu9ziBajj/ggojB/KkpI4pR54rGHoJEkz
Tz8+dmvN5CHoxdJ9JxKfC06SqsQTMzwVEgK6nCkKLVjPoJ4SGhscIEfDln0zXHN3
mW5P7e10A33x0FpWmK5wKVa3iqYgdfixmxYH61kIYU8xXFa0GkHLVAuhdDuTZi92
h3T9iiBS5rSHsZzGsvU6ht0+GcZpyQ3bPFXt4g/UyLTpx1Q1w4kjBhF8cCgCClj7
83tWajvS98hRNZXA6NxxBzF/QYvfW+zpXp/+cCVFmBxzN1L6EmO0kQkQUBk/Rh2K
gzVHHLQurSYlp1l2+5Lvr28726zeoI4RVQJR61ZhQ7Bs0NbwEXjF0Wra6nmKaecb
/OYxcqnX6/DzFJ3wfzBxYXFd4aj8F+qwP3Vw3EzO8+0GA3naN27EDoAfVH+o3j8h
IUCFCQRxhjnENQZ9yJVXrs3B7/4xVH904A2ka98BuQ3H0PWS9biVAxOL9xWa/Q7F
TdrZkV8UvAIMg2DVJ+cR+a6DejnyNHS0uWZIQAZkJ8laLh/Rv7X2ZoBfvo/Ru4Pp
ER5I6AccbkYqFaZjEOZ6hzmyiHYkWVhZSwKgLZ/1AR/SeUNB2SQ7uFnPGyKdjHNx
nvduYh79bWOfxiEZma7a4MHr3+2cw30ugoBrzXaK3kd/dp2zCmOk8SToxweTqUKq
GWryMF2AasKE0fBTyXMJGzo6rcetzAlRbKnw+878+s4KG6D5lg9ijZj3ZFuAWdLD
/tCdhBkHKpyPi558UjYWPQPpxmJQxjCiKrDmJeVjLhXj3TRvz3KUSyDnsdHdDtC1
jVdhu6ksHsSOt0zs5PpBna3sGM7qLlFsa0DmM13cAk+LE6GdPgQKRpxaYOklzXpW
VxaMJagJV8bu/xzNQeb+lV3vKg+MlIlplAT+Mwvh+ejkXOwrtD0THsqe3Mi0iMPi
BvWHyPFcn7yAQnuqm5SoWOT6BJ0YReFTdcag3MtLQUcQajONiQgoEAL0NPZ78eu4
Jtc/yy9oQ+EpdXBhYr9FZ4NhTzdtk46oW8uuLR5pClgsONVB0MWjBKHtpGwxlASy
Tx8UvAwKZis0J09aJNmHxNERTtjQHhm33CCxbOitL0NOBHITBGmR8nSZn1IiZYrk
o4WSKz4htMsxgF0paVAUsYH66ITKk+Vm0gATJ4OqeqUiTGj7xs4ttbZdDB972Idv
VXgAWTBRguxUdhRqyjrqEBLshbdzgPr29bGG7jOilCQUyTDsBT7FH6uvMnptZdJk
wpztFuYde/n1efUZUMc2eymOyeK8IpuGk37Lb1Zvs7ygovGknsh0bUsdjwEnAn3q
SwObah+vt5e8sSprsPmNLpwMjAJy6WWTPhmStkIAp2AlPFporqV7xO0/mcY+lJTQ
yYX6dfWzgtB+He+0uO2kiUN2mah/U04KdW54MFIra2HcJyziLJZMS4Y+m/d+4NWw
f5d66n0ZZscay4JHu6h5Fk/DwhgMbVaZAX1f2CvlIb4JtvSomtg2+fVNZvYWz1Tk
oXYtY/uOPwNZbvOtbwmzJHcDQNqt7r/l/dXbyxfaONxemjSEt77iXEmzG7ZIZYSG
32mGjvwLQxQmLyNQ9/HwIFnigURxAO8Z27eY232iVr9N5AqyuecZWRmEpy3KccDX
xWSCmQIigRc8JIsrDW7wM44b6ZsD6yvZQBbr9AE5sTAL2FhrurpBLCzCzNxDoXcp
Ru4BfM/I0HagygFNIDmUiuBG76FFIdHAKyiz6MKGWswGH4z6H69EQ/oO7Sq8CF2R
7BA75qhtZO/4hOgaqJIFmnuKdK3W5DREpZ3AvrA440aBfai5cBFVlaQgKsRc/AW5
5dAfTYM7QMUDg6q+wHFjACwyFPj3+geQ+WliDXFws7iLHf1UBQUaN+h03OCPULz8
sVlztf8TzYKuFU+pSl6rgaO+OMtXVjRfcABoST/g97uZ0hQnSYmOm+g4oJ8jyodY
phL9pkXSarnXeXtUr8prbFWtdO4AxEyYa9/f1PU96jwwNQ9QmSl4utWRhVnREVRl
bW7OEFW8nRaEOShPHhgx8kKWX8nXB/mxG0wu/EwURlx83WjkR8C6z4ffm0ODJ4T2
QK+WyOop+hmcT8k+KICoqusmJ2I+v9AM+YHv3ZlbR1NqeWSXxsgKPTNOIMcASV1c
rIc5RlhLAGKd35RT7x9TQ/fS8L0hCg4gcET0jCcA0euiCjJYHbb1mSfKdV5yQsZR
lbIO+WTlevgun5EIv+T/SXtp7wWfE02tURRbjZzMskXCAYgEo323y0WBFif+oEoO
5k+7e2d3S/iTTShwENGQiwgE+DpYkaopS84VD2i6p88F5bnz0Y7O2194lXVjTbjE
e1t1tNLpfaDDEyINhkCYPzTa7w1iBA2GtxSWJESMYqEo/WgCCjGNCiEM9VSF6jnU
hIx+0/IkvkYmcc1Keoh3WIGmrWD0DBP/A90F31SfonLybCP24PF9Aho5/PVTcDaP
7o2wu8BEeIOm1CwwPx2zdP4zTRr6bXMoChEXmjrQzSyD/mVSMhz9dg2t3PzQYqqI
rs5TC8wbdDAlMooMIj7l9gXwvDyrSoJ3PvpCzCD/FYocmHGAG/CQJ6xKbzfYYSvt
+lEj++XJkwz60KDMovvYW7s1jB0+ux1BOUL5O5T/5ooDWmc0vBEzaYpPuxWBi42G
wWe5z2mDwL0W9MmpybBzZs4RBqaHSvkoAaMcQqJE/WIME3wRwpxpgWAnWGsCml3m
AdP+rNP3EH2+0VFe2QsPPehtDXMq9vi98JL26Grd3O4JDl/Ny1p0zQR9FuarYYkz
G5Oob8dn1ayThK1OViKcO1cRUKYPG7NibdMS4wbO//Dl9CCKBkbLvXvX4sIeoebO
CN3H/a+CCd4I2Qg6CrkbSqFoOUEWFNE8YTHbaPIZ7I4E2NsBmUcM58yJwbpqfkzi
lJg9nvUwpKuzmah5EEGUEUJEx+vlAXt4uzpHbyd0d71FIDwMUyljQdeSOUJ8hr9b
K71SX+vIRTIjpK4VZOgjgmBT1U9izJqxkK89gv9mZW7QQCGtwPLSghVuz4YYF59g
5vLjda2Tc7TEppteP4rQ9eVopAEsZRjeWxKGFTeZe+srCUGCyoPhhvCEOGTH6FAr
t5bSutJpqAqQB/IMeVgH2a6JaDEYO10WlaHY/3NElKS4Sgo28SJh9sd7ZBhL0SIx
KoPfh6j23Q0QGTeuWOoqJGxAV78FoudLCC9UQD/UnhFWOUTe4uk5vrvmwXVgbub9
O7l+per8X3fSgifgdWW3hqua29/blOELjRRwQ8DvJ+TTlpnu1De0tahRK29FVdKh
lKwNAKB++5egbmNOdYhykhuaVNwgI10jV9/BNteSoacRK80cOw4DX3G72tU9dTn+
4jnJcnOGIPf2gzKanl85WsKX36S2LYpLwZjMmL8ZLn3HZm3A2OgM3oLKtRQZ+Hpc
DK9NVHi4nNNM2a19Chil1t397566h03urffwNXdDNJKcXuXwyq/AKBoP/M1Z8bun
WzYMP9pLLYijGZBMLPXHL436hd7Kf8NLTleqdOGtPaMIYk7RGlW4531rn/89OEYF
mSUleT7kuEZQGpEYWr/8tLk2LcVhjW5R7OD6LFFfJOYs31r2xD74dUoTqm+S8Ahz
xUwaISYA2GxELWER8/CTE3IVmX+0CQkFnu7PR1Y7uTpSPUeVVcuyFK7uMMub0ZWI
gBZ4xfdC7TZ1Liw4ekB5am0PBm6CQ2+aQJ5F98Te+pLpmgBgN67eVCAYiP9xXu0g
4JRwTcCemyAWFtqfFabNqA7SvIaAHPDwnI6LcYWdbOzr/HOin8vx4QmEUys1khYd
N53rPr4K7PVfOcL3M0CpWQzWXrVgJuRIPBr/uwGQyUTKR3nRrDoE2QnbnPoxJlYX
55J6PGyzGoElACzoOsNsGvjGZsLatHvDiYqVPHDtkaXWkaXsYtjvYlGq0onyQc9N
92GLNW70dL3fKs3c2Xgc1t7SOnA7BtI/SIDAMqBYpHPRnBkhRLwudOr1u9fDvYlH
9P/tTfS5c9SO/njBnnM50sAcUfg8AVFQup7Kl+kltkPlUIGtjP0/yepOFYtEqbEv
WISWmJijS148URK5yaE+2LMw2MLXnZraq9e88rJy5gEZ2wKXuddEt2JfT9QWTekD
T9WqvBYTRsnx8QCo59EA97m2WU/F/X1xhgCFXRxYfQ/5yZlIaBgo8g2kkWO9aqly
pw3mvcBms52DAazS85Zog+BDrvPTMRwfPHoxJo7fGusgrVPHuhYtOcJ4sEJOsr5+
AqJ5vkqRHGTDISel73nzO3LV0MCI9W5CJpXYwW4FW8VPxQj4KBqP+mLpMwNuM+MF
2zMD1anea5XTZiExQmrjO+JdccvvCI6An0+7KP/1WQ8d4tTfwK7EYrHZJ/vKN762
TWyq6p6f2iJuVzzvGoShvH7Nzq8A0NO6C38pWyKGPrnF6fGpEv0lKkEaefQFSU6w
Wnl7T5IZw8RqlJDb3I9bMF+K+SFP7YSDs6ZC5OZ1t+fgl3q2/BjhrOKw7rS7NMst
iOyEW2/C9R0NDVSWBRBLHnhuB2C25fThPz82llJcg3zsyDj31FEbT7Kaf81vFout
ytcWU6xr1qfmYRWUCvpeIFbOqnDGjKZa1XJSnSGCPEXjqDrg2DZZgI1XhEa2GM3G
Pqfz9KAt3xAbJNcUMsa+tnaGb7Dc/cUu0Ddr0iq9OcaunFYf4y1N8h2paB9UikjN
u2DKa5cLQcE7YZDvx8wvIFSleDEsHw3+J1jQ/VxcfKZI0OQcpYsxBndfuUvaTLFv
ztwYrQkK5mBwp+Fd0cx/O7HAviutxSvCJPcBMaD5+ZurPMm+V1hp9MqCJHvX0td1
u6pKCOp2LV8qd9zXayz8ct1Kg2VZsVb8uHPUdNpT+csOJnDKpP9fp3pOtMjNICkT
V1mlMmqpBlapf6lZYF6ChLWH5nfkWGla6phaqAE10gS1Dr4y5EmOlf9f7XK99nOM
nTPn8lkG7AN4RDk6mEs7D5sAgDSsfYjjELfr4K0Oa698aCsU4AMPc3zyPXDY5u+m
QwZchCCoGk1jQc7Ssnc9NvN2IoXTSINK8kZfXY/jf0PlM1hvMU/bnr5pa7iSGltm
jup1W7pC4RzoM7uYPUEaaLNbaG9AEVAFaI2f0GUBQe2mWgTMxaRBWJjuoUd8lm6l
2/cridnBN1iYvzuIZS7capCoYZIw4lMwclgOc19T9MQPlRrIHwRvC1cMYvQSp7cW
/dFr5d/6IczodT/RlxLTrKxnsVo9rW0/R9Wp6DIDbjOclD7akij908pCJ4LSVBlc
FGBUjM7bbMEmcXVGgagUZMM7cIiS0BZTwG+c8IsRfO9aT/Du+46qpoSsUZEb061F
2dSu99MxOj/ugJXXXm6JI5ryNaobtFmiRsAn3fgpABerX4+XdEjqQTedYfm/tb3a
1qr8FeiIvDA6z1A+xwmBWDR/RQF6HkVrgirSxB0zRPV+WKfDnABtI66upcH2QH/q
0D7FRUEYV8sW2OtiI/TwhutcVUzUqB6j1SPMeUqrR3x6/8RUqUnrqrU7I72E/28k
G7vv16hQAoYhMdCCRlmTBujWZ5DjWxDEZUvLi7KvZYg0dunJalWanQd6u4aB17cx
hD2b87F+rcuDrrnPdaYaiI/y/nRSkbwtruDmoIZwAxBh3Yylw6rv3LNAaZxF8wOp
iDgdknG890ti6WiXJ5PR+XWeR9yfbc9W1b0rNgpwAKZqs4Own6hwAFSVDmBrMBBO
TRR4wN90N3qoPlszmqtq6HtcbO6jaiqS8QQdv4a3+wbf1wPulyhkuX6wO7tv6mra
YL4uQIsm4HFWreql+OoyyKgSKScq0kESOD8sr9Fq1YetFyMEarnfkWxAVOOD0huF
Xob/VyLRwLUO9YBsBQXVbf0cxOMnG2VHVYT3vplCiVqOcurZC8p6+cPKxKrN5JtW
KSRqzNpAstF9IIuhDcMGpdY+an8h6HDmDoRWUMzetGKtIQwxGwTlJBQFOTBXeVCn
WhxGwjl3ZDf0GHuwvYogpKu302rjndSwfan8B088ZcU/j+8+uKaQMc+W8gdDkFgV
FG1eEdGICprphpZzaNnOceYsGviGDtUGnNyqlCBypuzBj+2EQRpW3tNNNAcftJt7
GVHbEu52XiNmGCv7Xv8stimtC5B1/mcLeNI7lwD8JA8A7uQP2YpmpBi/Ak+ovN1W
Ov/uZOmPG8wiaE4pciHNIcwjei2e1DmrP+RAM/LA1kO0/i7slShwoDipOF3qDV2G
boqkY3/BPDUE//hvZqV3svfCgH8+cOZVikPmPqM8XTkWPdiETFmmZ0bKKYs8q0Dj
3POvvEdXo1zH8+2zxh7juOjYZFBytbNkuE5yo7BL3epK55zhVJMeF0ACQGJh4fvJ
/Aembo6RoecEM8uzaX1X2SvljUteI4Mr936iiiQVodN+rkJD1kZ5QjLxwm2RYnj8
e4r6D0nCsbiUtSLBweRuOMoTPm9oamiGVM/QQT1aEiAsxJ22maKaIKJWoYgkbU/Q
hQgDX2LOkTmCb6ukWHy/uI9i56qLzCz5Nk46m+vSdg3Ha1fTPZ/yBdk3Hna+B9xQ
VQtHMxQ6hXtBS4ySYiUh14eMm4eIUd4ofKT957bByyapck497X91oJph8VoWwJ8t
0XX0Eff38hIe0IdVaH/P/GrHNjOI7BFMLyXOeM11qUVtOnK/5LRqVm4VcLhicztK
p2HEeMi21CdO76IAcijMazyOvcswFem90ajexxq95WmxD3nL4uy5/e/6NYOJ2F64
0lCmzYWbSeVPAxvQE4XdeHpcsEXYvi9x5rYgjZeKQrvOxkDmXsinNDgMtSdLZMww
CJuCYEFXTdxFNGn6lBHvNrt555gM3ddRc/jPfvpjSugCSgPgNHjvnWlehGmS+v3K
ES2/QBzJvrHZ3ePS9vxRy0qxYs4pG1bLs5j2c4PoqvKRIGaLXyLDB03+10thiw//
30sKWUsbfnbE+K/I+6lOmqxH9PAWhcT6FFYddXkxATDqAzrtOAm5GBYSVmS6cGNh
OVtdvgoSrM1uMPPdVO8IxhQeEwxWGwbFofoGxiez44VgJDI0thtsH1klyZEmbGB2
X0hbPzHH5ttAXpP6kyXae/z6SO2HdLhtcHfoV9mKLy7X5smH/MMHE6uxDRwXbpgH
Q2RU+beFlNZHMAaXP1Pj+hYgGflV4Tt2AGzN6ji+CdzpLEgcHZur5REbyK9cKdTc
LCTuWqyDoN3pJB6ozmAcN7kTBebzzbMG9VXSHLD4q1hwECbT7QtBTq6BYqlA1pwC
qTpc7hN4sb2OVuN+W6Lg/1EJHqG3PoZ70uIEtm4YFIHTAxMI0O5lDEWMM4uXA7au
2Ka0v3zMrAmRZAFK+hHlsrg/+ut2k/0PFx7mJFOojBeYA3AwLnDUVm5EGfbszG43
/kjUX/yVUbguVOXEHX30FomldnJVHsVOAdx4aVn6N9l2PVrje8ijXMNWn1/wkkSs
5dr0m87+XWJEfVTyGP1ckmBMdnf0qi42wIXDYSPugM8tv+Sq/5VITHHj0e6a+IJB
Ko+ZiAv6UD3NTWTobiBLLUiRw3RHzRTTLUbNmIeOfN26BcKpsGyWDXu6WF0BNoDv
0ctd7IXnAaHNc83e1n+yZ+IsXhhqrxLi80X3Tf3L+3+/6y40mIY13ygOxZ/s6WXs
SsQv5t1QzbRW2BPlKmrmQjS239LY4F2DCZldJKjAvRBLS7JK5YMWoj1c57k84okk
3Bq0xlxmoUfcJrhbkDA4pdin9plzZcBY8Gvut61sg8wcXYjX0QxKnHf3Cb+vHHfl
iduDMB9sfmrZG1GQQWY6s9eWW83etLqyX2nrC2b/XV8YFP+YhXCwYKTD68ZNiJvg
luor62SdoEsHG1Up37z1jDoCxHWK4MWcHJku8zEuGBCd0WQLarVhOvDV2NjOjIIH
bcObPXt5zB59sdO0nWTwmyiMQUFY7PMRe0WKA/vYyhD9sRghwf7jzodNV48+NVi7
6cPAMsfLlppnbF+GtPfwO6DTbVJil0p5sUnfc1E+hsHqH8/tiCUfv8tGjGcdGyQW
O7xVAkMQCqk+9EVWqAp/Nomg8nNvSFV43O40mjfYv5qwnrn5ByGWK5Jw8LI3Sjjj
Zv0kDJk0FMAPcWPftZnxRqp1LTNFsAk0XEbzsl0rjoCSo1Z8ymJ2e8FAbZj6sojH
My916K9ezJ/RgzhaUis7EPFtNuu/NmHcKTKp01yJZjkbtZxbp90pNs6Jot+XH5px
O+YJePymC5B80MWg2ImXKZttE41iMTj7vT6jc/1OxaYx23bemkA0Ab6LgF1rEBYH
F1hwTOGU/v4HIPj0vQzg6E/3uZB/PmylhyACbpwLqYg8rLMqeHHNBdxonjcI1c17
BG6OTNsVkBa2WhxLKPnXu0G6WntMQOwCdIwr2t33t8cUCe/d9xxWOFOR2PbEw9NF
afBi0M7P2Pu2bAhtE4yXQoR05FtwCJHzE0kcve8CuS1zG7Om6pMOumRqj63Q6nu1
CZU9WcNTEgQNXyglif5FiQFILBkJ0QR4crel/+uQjEnjyU0OJi+XY1DvDA5wbyej
gfY7tABX91Ny5RTW842O/NXEde8HI+i6anVsMHhN+gWZgJRXoBoraViJ7m/3cFxb
BkW4l0gPO1SjcMseA8VUmzNlVHjVPFOZwvFDqaidTz4D0OVdcwVqykRLb+r84pCs
dyNeui+9/OlWGipmJ++GR0gOM4eVGbzyWN5MLo84zqNXzAxEsFxQ+9nkYEcDriKK
Wr9I4Y3F572DNT74vj36Kd5vnxnei4Lmw7qgyA4h4+cSq01Lag1wHx+FQMoO2EYO
ZoucDWlKe04FJBQXDgN+GFWHXD3X5flrxcUDWzFL05aBex3wrKak756oCyZ63k9V
feQ0GoqRz+cdw34Iy4S2qolZnpOvsJI0pszolqII0p79EfkpnWAg6Jv8WInSsg2y
yD1hxBmD5ucg2adq7xJedqRapbwz45BRDmTPMS8wTAigLSJ4Bg0dP79g3UyNO9gg
xBuKkN0oB/xkn3NwwiZZrFO2KTtTSwM9XrmrVQINAgZJyGZFNnbwSQ8HoLNZs2TZ
diPTiYE62fZKcgN6H80ZCSjA25r4nhvV8ByVFesWM/kClSvRjaxnGQDdYCXCa2lo
wnX1bqUVUMF7xBLp6ewtJZgTIXmeEVK4da+g3dcE6HE8y1v2OVNOygKZL0YD808U
2iTPxPa4VmXes1MbT8LuGxIinW90kLvXxL22Iyn8tM5QA+NJaLjg7IbXFNlec1xw
GfKUCwbnCLtS81TqWQlcEdPcoqjLc1bJEw5ve3+bAP4seSSZzHnj1y1iZpvGOHxi
inZXb1aNTiZ45SuVaCuccI5Vw5YXTJW3972y5RjygfxC3tU2GtGHmkOHzc107fYX
zWLEAOLC2dH2ffpbS8u1Bf5ckM8WM8piSMra3qy4U2BBZPyddwi9yQlaznC2PkyI
eebDH4xU6hhHQGS6WRl7ZBvDkVNAC4WvGyQsteuKJVjRmaJqqwMhGgixcRecBC6u
Zq4MlC7E3iDzGnhAC/P1N68YjlgfUSUZ/nhOsNT2d4pbjcmaZxMXeGsrpHDdvyS8
tDl10CFWrJchUQiV9D7fzrybL/SlNR0thh1ChOZwbRT4BRbDCZRk0fOBboD6rgkN
XJUcRDmGRYzo7VVu0hiPI6hdFYsfOQ7plNmRaCj3YPd4MNCBnJ1+PbdnZgqHyLrs
MRnVPbJaoPjqcqQ0HgN1D7Gl2JtlWYxCv3l90R5lCcfEwBv+vPAb/u87u/1Lqb4D
twMod1+ciIw6BP0VB2QL0NEzSjTHbIMqPU9d2bHjHdZQEMV9ikjurZQ0CgYTkTrS
ZmgRfHjOEkpBaIHpzxNKK6PhF3NBkvRlTipmMklOtFaKKEMyvHQZsTl7Y+x081rK
PTYxXWk/ZxIV+AXPmg+rKEzM65VJahT51Gscz8lQMXOVeiM77cbgL4dZDkVhQ5lf
6c2/OVtJQmB6XJ+zNsgfncX5adZBBLwaIshgs2MsgGodDf4SvMyGV+8YjBk4/wio
K1PgFIukuzHvbMlgCXJumQZ08DiBznXMegEDK1WVBlf0lARv4Y8ODkLvnp4N8uAN
dZZCL5dZg34pC+iXSrtUG3YgDQQGCvIjrQyGTLbi2xrEmKeOK78NAfJgL2Ec2uuo
MYK8DVYvgk2Td/AVqQa/k/6iyxa9APuOvt76ThpDMS1jLwBy6F+SL+aCxn9qTums
9H3wGDNrozC3F+ZtpMb0DgjtHd3Iqo9ag4i5lwqVc0Dy1tGI9a3lryi2aktyZamd
uP3p4afH25etuXoYgdBTjIVsGwV0kHDfYGg3FtfNtJsXKXg4getW5czT09TXrrJL
vPeWbYaMX57y3TqfJFIHgCdx8FT+q++6QRXx4f26DWa6gGC+7e0DjBuCI+hUegQk
90nGS76RDo9mQ+Ul9VQ/G2XXCAjnTKQR7FPsrMFXTnlxxOmoZgpvsOjGq8DX2P1f
CwddwkEVO/8Zh+LZSCuOHP+5iz8pOh0fecq4A91TRcVLPk45bBnMp7ZMpEDZDAMK
2xTybr8VX4QduZP3JPPp+2fX2d1nqzgyXpBwLzGO/nEU/5cyWID+SOOOEyc7fe9d
wiKlcEZFo1Hlyrk/jx4yCRkAcEHvGDWwc6kgUQ0pzbSm2ZNfQW4SoPQMqjVILiAF
+bWbgEVzlGe0vzYvZTKGeHtOUTK5G5l6Nv26Kz+zXf5gEuh9/mbM0S20OG8pJfGZ
lv/xB3ef6Lmr4rTTG33YuHK0ozisapeD3OF8HhLfUWgVLNyIhhzkGxAkP6IS9CW0
dsTFH5ErRlDcgl1ZzWwuH8N+RV+m2aENjGIATDB3ekogEuhWdUYC6M35t0OxZ+XX
xBUod7OoMN48uibwJXIKnJoLJzsqy1DzNZaTMyEIvoQk5IPlrOxNYSDja7H1ydUE
523CZR09VDv+Y97crsEG96FTu3+BiuCcI384Lh9ptxzv2VZjL3hDfb1pzmBSOx/B
SDWY06hK4EBZyYPQ1Kd3fqgsaItdfzrM7i5ENHDc9CsJ2hbLyTjiMiE6rQrLTjCC
Zcq8+8TylTp940v1VUZogYaBvbUWRjPcE30HxTABufU47DmhbDUIY4q8Ahu3j4YY
iVymOQ2OVjWhAa6foOwrSAIybMbGTx0CB12hLimLk7Mlx/JcfnyL8cIZdUsXbBNr
V3JelhFPAdtaxOxv2CdkJKcaY9O7tRvYWIic47kt7KUkrA83YeP13B0iqA3tw6/c
uGZgTIGU8Uu1npuKEEwB2aZq17vrv2ekZIJksgdR/Rg5MxfXand/R0+5/YQgDbI3
PXT228rTRENgaA4aCyr6CnsAi11U0nz0sSbd23idYQO3HiGS8SUVbthDTP9BpliZ
BdjLq8ekDf/RgmBuDmxzUqkRsM5X4K1meg+uz3EapnVFq0glKVHoEb5a84cfwA+N
YrZnV3+pNW3RBaMUbzOVZBBpYWbOA2eoS3DWoLZtvproiqqS+AXEO5vv+lnGStFD
cZkPRIFFisqbn969pzkpyDYTH+qr/UMOrehmlMoSFrI0zZWT0OXQtJg/jcwybD5f
l+WiTbJGJDcLxPuRZTWa6oFU5fcxFjXQlN1YUjJQOuvj+VWYqpv12DuAznCFdEAM
l5ItJWP7ZUCafKgUf0MAbL9P+xtydlsIfZ+WPC8s0k5kNjudsLU1YqR69tn7gQPr
KvJ/K9sLUEBI0fQi0zw3vCiSuCy2TKHi/WGsmp+jYq6+M3XWrie8DRGKGWDcaEDB
nBMLg+BJKczSwqMpfHhHgFfzK2sr7TJVKspaA/GKgb5mRkQ9fF7InZldkAC9dmCh
n/gcnjDhDwI7n0vfKcBakpauJGM0+/zUFcy5hcFEZzrUVwe0Ps2Ugw/M7QRiTe36
QLPn/pzE6rv7y4/HyRq6ZcsQ/hx6keFAc6cwhXJGQx8iNfftHPXhxflL6vTqyxtn
pfssOi8OYKOZSH95v1Qq0WPg+C4e9CVVL3d7DPWQv1t0WFB6uefX5dtr/u0mROGt
PdU/ofsqrB2uKI4a65BAzYhkV/uENxNmc3HmyXjKjuiaSow2WJBrqByD88gH3Rn4
XjXfNVEJTNA6RsOiHMYpJokU/QIuRj6/BPX6+oi4ldk0MnivIoNDgiTfznEHzDCn
jcwiJOopSxmHFWxAyICtqaZsMaZAWhh6ROgJ6V69cj6xitnnf8ABNdF74nwLx4Jc
BofKPIII28Y0gB6fexn8Qr7il5VefWQKzKrUilW3vyXHJnKeIqSjCZLRHmm9RLCi
f+yECiQ8v08Fd8cQzakBfgGILGFjhl4EKL1lX9RvS48/+L23UqRJXf3HQgn8oLml
nydhdGDOX2RRXvBYtubIyblpKsiI0GYO7W9lED9rBzVfVjjVtyrTSuSXDTXiNdt5
G1IvNamr9tF1rU83VvUWMAGJjfFWYg3l1POxvhzQQeUqdKx4trgNFxmEt3IEdXCe
RTuWXSpUtAnDIap9jjBjGyumeUZgY8UqsJhCLLo/pyzIRV1ppYbo+NK9mCgsQVIK
q3xeQFB0QFeAdTlWkVIESYlNEogcUXdSHNvn6e368tn371LLE91ZqZJSu9PR4NhI
kFtr/rreLmxlWF+QIrJCNzgaDo+BK7LgroLU4Ebcj5PIYuLul4l9Y8MFTTSZElei
mPc20z+X5wxfuhQQIiFSd9T4ziFFf6nyFNsi6YMP1SZA6ztZSPouE/77sdYoSXC4
2WDY4lpQ+aB7f6cgWACR1GTkLJDJOyFVDNw53H+MwW/exIqR/dyx/6bkoud/LouO
6HweCFtjGP6Mnv+GEeDqvhbNAQmCC20cL9COmalC/e2D4vLkwrK5t1HPu/BJoYyy
70hDkWEEJ7oTiwW4z99fRLiI56bo6eFKSgtowrhtLlwfx41jjIpCL0dalCGaZNna
jBPnTE3enZBD76eT8w0f2sseWXaIWBnnhhljAQSh6WT/MQIrQJzHmC4pzevsOy4G
ZJ+a9QQzKKxt1ZzTy0Iu0HZ5IDR3pTuEjDquGyuONWGuud2i02jyVkFy9lWLnjW5
fG6v/booUbjaiBfxoc7Q6UUNmYV53HwFxTabc0NMfB6MhwbnLGImlt5Dy7SoSEFR
qS8K9kJDLus/W2zLvoW60IxL293748qEn7A4h5yQwp7QRziA2sREE24RPCqnCkf0
uN+7NH7RD36ftwSrMUIrPuduz1wcinZkDA62DBUNaXxdINw0DBanD/bO/nTpHawL
HpmRLQ3ogKpyGa4oJJErXzdT98qwtp47ApcpMKTaaPnJd+tU73WlAfTttwnwqs0F
Gt89dnhG1HW5+FQGue7qrbq2u3VIm3c8zHjsQgbPTXy0psFGERgaQOyVt2MO7l0q
4s2/z08Horxj4hiUL0kSkyeRlSwaeIyaoMTixo9zDLmYnWzUDv8BhXqH26BqFFew
IHnMiDmS/SkkSwYBIaqXLg9R4so5Z0dpP/eZtNSItWArft/XKrqdZE5U+5j4S7R6
XcxrSsFmdenm1yo2I6y36U8a6N0Bnwa8v9x2WuuWnuyjT3syz5XbpS30lp71D+sY
AG9H5FOkj6vwDJn4rPpOUV1BIYZRfNr6fzLOHe3h83foid0KjEFbWMhYDrCkodpN
KM3OZe28K58pU5Q43JNxBIVmHyn1NvU6XCLiIzHlkwnxDq3VyJz/hrJFMtw77Brt
qCGn6An/lCQ5rGlDM1a00blUA5VjPjrNiKZZBWHyzZYfOQ5vzu5tu+SGOwudOEeI
iFf04Tjh2H1qDFdJlV/7ggoJOLIc5FAbAo0jns2RlcuLpKRNBRINmywqEwqEjcg7
oaop9JhoAAzSxVPuZRt9/0NSwR5kVT8NdOLItz2a7qBG7XHOAfHp7GTnOMz9c8ID
BJbjdLxTfybco0Gf/YF8laZKltkEoB+fx20yBXV/Q3ehCfKf6nzEw96Tl2quV+ze
UWXLHtItDNx2XlV3d5F//hk4+wRl7b5jzzd3glNxCZtfZTkQRnksYqVmxOsnC4cj
waP3MC7thr9pgl8aLAOPrQc63lXS7xXTo5N1RBw0yHOUQrHLMTTYBwUm4PWLBSOY
6xSXf6N4Hina1PkTEzNzc7e5woSGQvheSvwi2hK/CJrO9nyHhI2Cr8iQUunQd+Di
9bQI236fibGJL2NWvNM26tQhZLPqvxHbzu4YhCm8KuPrMt4jvVh/1wVcqdsdnhIB
ofFOoaJJdpBs3wiCg0fCb5QV89ViIulfRO6VmvZk4SGBRyVo21B8zPcabRnn/w8I
NpB3UyAvUbYsAx4gDAf21TLrP/hix3t0LXORdpoHntAv+2TMHbxKxPrfBym5uLOJ
cwqindnw6zNGQgU9gh84CPjErSORHTbrKhXvTn2boTiWse7NFBbp1MvRMT3MW2UF
u/CzPqhmGU6NS+xXJiLLt5zzgtU/ZG2OIk0QNVM3FO2CV3ZbnSvF62XpZqcWdipn
ZTZ/UC54CvGO0YmmJ3b13LQxKdG8CSTjcHoqDXspuJcr9byhOdBglWt2FA2CprSb
UQUXdVHxtGSYeEoMD8ig6KsVoT7MJqJ7hEe9OOh11KJzeydN9pzhQjREegFEO+tX
nn3adUCNN+UKuei2hrguEaxpUk1Y/J7IpCa+H1BcHcYeZ6sdIWzgWgeU2oG0E8va
QrjdnYX6qE9Q/DMLq8FF6a9+bYILggyp2LrWca2o+FlFsv5rG6Lxsm4ElYGy4lcp
yu333G2J6WnJII/1QGIteMwAn8iTZYJ/5Iv5mlsI0VkKTMMxFtIz2zugtYdlH2TY
v80JcwUmtIzx6aaI4t/LuJ+I9hHWu4vMrgfQE7AXpFE2Ts7QmgfJTw0QZ4A4DxbC
gqCfdaDjizRz3foZIKBIFhl9x1ov1CAGOuAWIrnl9AoYYTE3zfL3pzxzAt8qm9ay
ysl6lGjhF1kfPgddAHssaK+0dIEcp6CRDnktMvkoMizFzypequj8hykY+VXqG5nn
sgkVgwxzw1WNb4sSLPhC+NKBVXdS6xTIEugQAtHzuDbs+mlJ4Ske1+hvrdgVJ5Rt
oMlHnh5bIDLfogFHSASbum54MvC401UthTbW5NbWHLesOg1koY+vveLHPJIxIXVJ
Dfn1hcp6RrM8rli1LTRcrqPtdAZOB1s4We7TzpXdf/BSJ4ZGXvBsNFtn8YxXAgcM
irlazJ5HLSnsY/wAxhJ2OQZPxCWuGvs1RLBv6LHiUtaVM9qHHbdUnAV31+dyNuYw
1QcqKto+cNG6KoVZH/1GCedzqHj4Pe6r91+pQ5+rONmxagAkiS7jvD9vJ4IjZNqB
ZkUEEpFvVB1BlkGVB26geuthv1eF8pI4gtWisuSwy6GrQI2JlLw/wwUMW7YB04Ix
qZspoW7/T9JbaicxZPFznNoSlp5+29yBvDhS/2qre2zz7yV/fVvPYaIjDibsf/C/
7EKS1ovAgL3KW+cDC3UkPJuegr6ce0AcapBEtOuR1ElRlh+AkgpgOVhFcW6DsQu/
9sAQX2lOTS3Uc4ZKcku3XIr0ZL6NuzPkC+z8eNqVjnGrv4rPjBDs8Qi5W0k3pU2+
BUNeaqYwGsi2o8lf820bU+bpyugA33QKagit1Zlwlbi+jydiys9Q7Do4XOnd1ImI
NRdOTQdh6Rzyn3HnVB7gdwZMh99BUUl1DBqdyAkhVX90y6rbZnvSm94GjDEOq3HS
UJVByBoxWQm+MTc7IozQjfVZtEKwBMzML1iu+oD+zggENdFHc7wyCNcfhbmtWxnB
1GfrHhZIzybVCPRTX8cGdhYIbpyYAcNpqhkDu92y9xOtJOEOU5DBT+Sc58XDTPNF
bHOOdczQoUWsGZ0nDkT0EzenVe1Qk52tW3YfpIaTzVdBexI5/6C3KRgBHeyWsgIJ
eWeYBVx2XGhQ80VQ+CHyx9M3K0OngtaUftR765dguYfA27iLnhBNVV7ZYXHsBaAr
fce1Qj5bma1TfgU7wlCdBCImLORmnOp7R9Wvrrbf8EOaNDJls3xn+hyx/gRBQ0Mr
Re84BxXflg/5sZG2joH7qLy3j9bjiP3pD2SGykO5AUQoNlZXfouOKJmZcypxHjMm
BGxxev0gUw7iPDhj3+bZLaqfSzBavS1gkTtlfinnOKFyyfMK6gcwQwgGYFGR6MiU
Ago6w+/Z3nPS+CGhGuXXPnAQ6DQg0HitH9mxZedAN6XNPb0ppK92wc88l3uMshME
JGOmc8oQmJg6Obl8O4nMGNghOwNBSd07h5VTIjIomcgOI9BSbAb143Cv06v2N8Au
13BqCe389QmMfsCYqqMJos/0JGrN+2h6dWwRTi8Y/nrA0ERE7XLD0WS5ozZX9uf/
0PgX4SCND6uOVNF/sUTrnP01guYg3VVn8SpLzrtK7wWYMfXWUcVJh5XBlOGja+ff
9JhOXQBekemBF/EnRhpGCzYzdp+HrcH+hP8PC+gOTNZjk9nCfoNbTuQRX7GT9TOp
gCpKJJMz/hhqQTGFskaa00RVgr10vbE0ikyxvGluII01VhZYV+Dkev60rcCSNp+d
MHUexNwu3vAiramlNdixkCKX1u57lUy34wZ5MmTbBhkcFG7+qK5jGO5yLarnM+3A
eNtACkMVOPJ9fRjFWb5JP4qBvfqAiTGZKPnh3fqTTF+IgNNAfKLgtpav+wWNCJX2
8R2Qg54uUW+9YngO1Vm0CAc97NG+asD/FgiFiPWb5cPBUbpct+fwOBjy/cKljMO5
5AuT5CmpI8ymqhcL0+9hXwMYuowq9p57Pbn9OrDFvYSDpqeQL0gnSqGFBJ5S4cDA
433PRA1ApqD7FEJctuw3Kuy8wyC5GgdCVUytSerM38BaIcZkJPCBnKNMpaz5KRAl
4fK7Us2S4/P5r7Yp03dcDDUcqAI6uGsGH8MjZUHSI8ek/giKl4l+PTn5c17gYZGu
YCfMzCwL//BGjy2HSVd7G1XfGRa9kyyXzJnCm8pcuBt9IOEjlaqOmJxzeyEwkpHl
Cns1Sq+ZqWuKYiHtu1WSOtxVSyHPnf0HPqFPSzhJc+udsudurXsCbFCbjwomb7FP
UKn+iJKvTgjjaZrctqdVjSu792czzIPP9gnwJ7nLYK8mfqT8nawVNHPTzbNroh2B
0osauox4lFOjzfl32XEkbXtg4lNIE1o10qd23JPgH9hhqKollH7DH7eTN+pH7raC
X0XkFeMhW0P+zwhph3liyNiwxCI92zM6w0IpUwbJLEZ1LDVEueejzyWviZV30WsJ
Xlkz6YzLQA01huRgTE1ZtccFIf+Eisiw8nlOnU8LkJEifQAAoh5d3NWRmJgpgAPJ
et2v1jGuV6kogzGsR2tFfTApryu8cqQH/7nXxYkknOCBut7zLNpOnKgoiScxDn5P
3xRFNgBDav580tArylZVXoKoETjZiEIe7dflibJl0nALqRZQ/aqVtaZYJR3Uy+aJ
E+4bdsAkbjl0+OdjRLmAtlJw7JhThajVYed/OD3UjtJ7V7W8fxGXoMEfDjSut5Rb
ov/ff4j+EnSR1IjXySxrYdyyr756/ZMOuSnGGtRSuNFZYNXq187Ws07V0jJ4Otqq
cN1zCKDM38Ep/bcptBDAejkvDjQoyGp2swXxt1ommN+xXdpj6kAseEh/JEbkmzW7
R3AMB/4eGdjmIjIVUsItcxhLzD6UhZXYAHKl2xzXchcahOWxIfMVSObti4K6gO7s
9jfKbaG1B8B6xGRfk57on+UC5qXdeQn3qnr+ev+6y+J/XYo3lt2K1yBjjpS+zZTq
f+3Sv/7zVHmcgnNK/6tRv/41AFDiNHv7TwSI+tFAdMha2+a3ZxQv4Czh9c/FAIDk
8m5WUqsf9mxq8ELGawDHH6us+OXGroAJk/EDA3RWa9TPlivBH6Cp9CxmMrnraI42
KYtC5/IaHAeup+hNWkIpuj/wlhrRV3g0rej/GQVLolZQxZU5UvKwJcfNmDRwet4Z
lb1JpMz0hslMe8Av1IL9PCPHG99pnULgQjx8H06ExH7fCYCBMqrl3sA75VPke/a/
i0noAm8nZdaj0xHmoVxpnRGLx39yqTygi+JWX65FNEv5qrpsvR41OoGOdR35p+9R
OraINoErp9VKwZlNDJfTQwBBU+Trn7AagbvpI1vwfjDYL8DuiUjnEQf43xL559ok
8rmkB3PZunr1OB7Wdg+6DND7H6m9dHNPaWxbxs86/wYIezI+k5Xfh3rw5682OCNK
BFjEJX/+ejUa8fiUfvquRJGtTiZojW6z7+QpLdUfbLmS49LstMlq8m3Jc06SoLyp
VEDJ6JWtwvqd7mhq31eYeSCJNpN2Fz/a40ykUZjfGz6OlrxBAxXVAaNW72HgNESY
+/wMe9ExbaG33aIlul1oAFzEK5KXnXvstt2UQ89pauAaGLcFIVhYzCKA6CeXyQdv
rDe4Wr3tut7fHbwWBTY5eFQoB4O9uaO24QKM2/QQcQxiRTRVUexGibN0qjuLciTb
QYy1CttW3OsojNleJJM+YjpatCRQ/jr/DizE1COuEf0kd/435+c65HGporfpsSpX
DDsdynN/FeNakrjEfjO/IC7PnZfMnI2NIEF0CqvD3bqBnv4mGuIYD0Xbt61c/t1/
HxqimHlnU8e1lem/bwu0i7tlFowckB67XaWocuB9Yq6yXq9BCYvpPIjNPjMhyTiu
bJLciK5dyuPI4avbIO0AYt4PIvznvif3LqPMyKDNAhiM10gJiOuO6KujqwxaDrZd
6MAwC3FFRHjbFjvQPVLJAZWkotdM53cTRPGrOklvpTd0HoCu9u8LSCcTmLi+qawW
T0OWrUieX9SYH/5wNOZ77QH2ZR5DjVpNfQCHkiH+s7jmJpCukwJ5TxLmoj4F+hAc
iUQcQ3VP/DEeuMg+wMGBUVAGM7mJmFrpCdWUhgxtgj/TsaRwX8nMl59gNf30I7dK
ol8hGWmTaTx8R0Vj5/vQAvSzMvPXlsjopzPL6qOr2cNyXcqeJ5acEmu9JuqJ7b0A
I03eFxVvKzVEHosq+NBh5pqjZc09CAExuaKaCFZQWzG5q8q74oQOOWeg+hgBY+iE
u+LWurV7x8I4AKOvKeux9X5of0KVEdkA8Bn2Xs0aJISo1r6cz80XodCezbSq/pI+
8Fscsky6ApLUcxIiZm9++S36ZAp4EqonmEgVYx1JGihWJWlO2zLZn9Qt9Rr22pbr
DF+lCSAHjCkpYOv4mktaNxJwCbQZ0FR7jZr9+MvqxeUQuZb0KB3+yhKe6f18hc9u
gBOJl7aWjbZOu/281ekEr8nBN5iNrF1aOKjwKAYdMjsEbu6LJ5+TdaHusFMZiaNe
B9UhjrNUSEinPIhyAv2xioNxDcyIwzDIYJ60371RavGsVSrIY1dUEIfuDl2W4oat
4npfMWl5RVFHQmfxOX87npv7PWK3LnXpOQCkln2g+4fp9ryLz31SjNtilaEsXzB3
petMYUC9AXWX133hx3JwwHKOhZOjzzjrNmbnc6iolFgsycjUGgWSAFTk4ZX0C++6
ihwOt/38VEyPrvkNtnjJ6gzT4SvYaWdjJDTr+Uy6De76lB9pO1pvQvv05agSLRRV
72jsbCPxmbn8rktVUwyt0IzcDu4GVP9ugsBmZ1RdaSSa4QZVoLE8RLyrL8WbF0sU
jFvPVHCuWB96/QvcCFmwWcPAf8jOj6wwo6eIlNtESvEN5ZBIG0Bd2y5kMgpDCnyw
kSzoMcRQIj4UeICw0VKVnl5W1ULC7CGQ8OxbmHLBrwC1hEjqyr6oPSeOd7TmVh5d
D99vYKsG93Gl6eomOJ9YWeNu4iu0fh3WVpjvbjmOAE7CQI4qZnGY67SBxOJjCa9K
7j8tLaFxN8sytzVfmnfvR9ch0Uktvvkuij44OBqEJHj0BP4tZLZp+lVDfVdKXjwq
nMibJptxoj3Ob/v8pdS4AOFj1wKY6hLoO7vIoDZkEl4QwE/90b7BPmk7cma0WAbe
CqL2GfoXax8DMav7gBjqmdkWFwk2d1XmDV4mQz8OfYtMXA3xKSZ3L2BSOfAHHzBU
yw5T1pfhbXLOunlfYtL4bEGDkZLKPVssPGXoptC6jXvfBxaPMXj8kzencaA9SwKh
Bh2yNnLjads87fQ7noo9k1Je21ofGytqhKkIUboizdRy9cGyDUs4YOBT7awHPDPO
ammfHH540mzzi+QVdfDcwv2097jxjNwBbFML265ZVtDQXxaz2Vlw6y+cuT+vSCiV
e7Lg4UGNXjeK3W42bmQP9/5R65GXJyoOGzk2K0vRw3q14FAs00fBCaeO6tq4WZzm
nzHMUxLHMSV5u28gSxQto5iEjKIG6r1/BI+OvnyzEsNl6fBMcjScpVtiWLiQJrMV
vOGWbfMPXLbGi3/z2ORJE5QT5VyRozl/gmqwCcWYotab6qbGBVAbpah8N7i75qCu
AKpu0y4GLh5J8vn7L2Pe6jwchy7ITQDU1FbdwthEe8xcCgWRiZ/Ye9hGhucoc0Hg
ySrwVUsK6YOpr+yuA4ZfxCwO5xCxDPQkVv7Ke/S9u/GNDqCUpwpIJHqeZdw0/eOc
4lX3KFE4vvirNMQTtB7LDpdv4J0Vjx1eNuPDjDlFVr+FLSiQgv8iF4PS+T3iw6tE
qNp/ruzUSuCrfYJv3ozktPf1qTYuLRluKKZWiyrTirJ48Gc9mB6iLuKOx7T/92Lr
EZDHD/qbVBALZ4gwS9g1g7zPfgz34ojfOuwxacv/5bpZvxRqHNdZZzp/wI3Zs7BC
5cuGhjjs16UfdwJ8x6UAh6csbTWj2soJ12pQAjmfTjC74fe6gMtmOwDfZ29xDu1Z
s+DBW/kNku3BAEtDbC9UEmMHGfwgITcF/LINWjQCppZdEe4CKUf+L9u9awr7/hgR
Fy7IwDFwiAFMGnQSTVEEHnYl2n8ZXCrQoDB38XoLBS0dpBJtxCxhvHi/g97nq5mN
Pv4aig5AOYggbdzW/BGV7DcI5ZzbItA3KrPzuEYZ8T65Zos1FHdiQLiXqNurdy8A
dobdbSrwbXyjjCKZSDPCdWcEBysRBHD8FdQYpHeyRmh52wViZL+KfEI35UxqQAHq
qPZdD1hp+h+TStEzbQGhgnJFpP+9eAvdqa8sycFhJfoXkV79CD5O79KcZQIl2YRI
aYR8u/kD48Z+uPJ17e4DbWk4JRpl0NO6Q5Y//4hf234gkaiupCDIiemg7kZfU29D
vcT1Agnj5bSyLdrxjXSRdSopOh+CYcisAdtQCtNIOQAOP8m0n1HlAubaFb33doJJ
XxNlyVznK6mbt8C5ikCaf7fUSkIQZEF+0ulPxADQ8YmtFgDRCnJZms7BtF9glaLN
Zf9+daIKA1ZhrZBlB564w2lMJGPVq/xXzoz/pGDK1s8brZU0Jear3wwPFT2rIQjk
1gEz3wT3vec+JUirKrum+rPSCt5v+a4F0Au2oJB5B7AmoneaXp84fbY9pBykvtNw
KeIfklCv4IcTWSHI7RgmVlJSsiqSKQAXjHuFMG6tqqZH4IJ3D3sPi8RTMyYZ9RGm
hAPMXS6XOBny0v91SWkcC4rypd7KZmfqRcIv6JbSHyxbyxAVL+SZ1+n1rMXX25jr
7+IEft9JhayVewYTuXlVEZT/7Kcyqn9Om+8gSZMfzLPgFlMnrl1CaoijmCHDIosa
XMD2UDYwpbMQt4ciTR5cucz+cv9QR9+vuX8mdhHR8dF5brdOfGWOdCuPmctFDOmQ
bTC36DtqQkSLXVVKyNrSvvxrhqqzEF4XBLVuDw9qF4F95ItIw7ZXkF584sFWe8LY
6mEiHhkEdPkJ5IvJN0lFvyRxpQinbs6i0yMh+e+6/sPAKgHZ4Xm98oQT/8dtvRUY
gCXk9vx9mPpQO0V1NM3bN/yDh6YSMiKzbJaVHzEMCVdGPwrQJfTl6T8s0SiA38By
YOWdFROc9qe/ahm/t2EcbKpPypzgVzc9ycuRPEfWa/lVpAPWZnWe8OFhr9XF89WE
QXDK3T+dK0hbi/F6blADMS8SVdUBUGN6sFnElpFMhjfVm9ffoaOC0D8DVI+zMVoU
BHW+RFeUaAXUAunx6c0yIz3SyzyICSfDbN+rjFgkhqlvRwF3u93gDkdCffcIlvQN
v6qyyyD6KHXOHHpLLsRU2PGRzLaG5UxxRpgmvRlYIfCoX6zblUCVV78oE0569Yz2
85eht9q5Fhjh98Z5F/pnn21rIVQG/otMjVxWGOdR5Yzb/3cAsS5HItxk3pyrVqbO
4tojgIc4aWVvqEQ/8NRaZ+6vUJ0ULtVyTbc63Xc63+4DTLycDv4+UUyVZLurpaoh
8p+B6G6YHXm8wkmjlLLvBhA9vW7QBoTf2yX4jSjmFQC/2fuAoCLI7pdE+CibdCcZ
7iT6/ErwIEKDLSYG3LLuOHudMd2Tmd0VVIhye+RHg3Zq7TsK8xKoxQjs3PHnekeT
UoFtLks495l5sbZ3Jmuu7tPmpatWEeSZN7+YP1CEhioy3+hJ6i1m4k6eATe3pbPj
yOxH5DHNT4PosnEyMfJBRiinqU5SpBQPdyTeDHUXmO71Q1i7x2fDltjrGsFi2mrD
y5xv5XxS+jQLJTl0Y8PSwyDBpOk5G68iUks1OtwSKEEq5WFhtVBcx70eL2UONOyh
hcmNqIKk8VJD9S5LsNSGMBMCqblPeQ8rZSPfeZkVhF5ck2l6i6uot7+l5Cje2KDS
UOWQz7gMdMcpO4n23c4wI/1zn5RRvS/gxzMf4w2Yy+r+FKTnwTbAnaA2u2GD7sxf
1PV7bkjqSxsvBzL7FQHVODIocTpda6iue6Ydc71d5z5adhZQie2oP2QnE9xypaHV
oIo3bbvRJKdnc9BraZOcqH1JyaXbnlKQ0l02LUJlQFgZdlckdjIkTSkvV46wD4BQ
HokhE/ssoDiPZa7jxMsHSd6Zo24bsAVDsVZVoKvGcZvtnwkkkJsOMxo6+4/zO3LJ
gV0STJFwLmGB1/F031D4FE76Wkc+u3wngMo0uqBqq6FXe2fKb8sZYxCABdputKLT
qLygYTKHy6WzYSIZ31Dn/8XaNhFMJuXExS0gSs/0Str1qVXcM7W0Wscl2By1tiv2
dbWFOwcJbaOedyaPqJOr39pHi9brRvOe6RIDj8dz8E8R2bsbzILwIZsnPC3zlGfd
GeP9unR0Oli67UkF4lnpJR0VY9IJ9L91UjOp7xCAwSPdxtsVHmLg15NDLa00B7ki
QZD0INwQW/2x+CUIiwnwZcxVbdYboRW02oKeigzONraSNY1BY2NwdXlS+LS/MR0J
dp0lAHHnAY1LF3IeTVI/vDcbe1fftY2oQn6/oRm9btb2DoX/G+Toru5B6qCS78Ld
LcU/+blsYK7c0J5gMAQjfTF2A4Z24WxLdatFCVt5/xSslGdL96t8305Q5z7PTxy7
6hr1bvrKUYzcPONVNGWqQ7HxRFIUEIY6utmjl5X3mc0hssDd+pL3iK9EsFGMlC3J
0Vzfe6V0YaL1KzCtfu1gWeZNJkfcgxTiG3GRhw3Rn+pe4EEU2PShCtWgb4RkLi76
c9nzuWX7ro8yJMd3G0oB15yFuACjQKbVtD2melxKzzQt8Amsm8gWohaH16B6CzMN
3YwkYWkXkdLRKjSgdxKJZvOyqR35jJcwH49eJ5Tp6vZCb1bLUfADrZPMn6NnTMqy
KB7Jl5dtWrCSYhYx3vjJSVjIrv2VM3X+hcgjKFx+y1KAv3ZI9Rr7NhrMHCMX7M1D
juNYGG2H9Adc2Ig790KkZUbUn0UQAGOX5Ot358OG1L4fnBCtNqTGecnDwUN5WEa0
cvgTxSjkxAnI0rq4A+doz02ZaniRj4fp2CQILtYXM6vDEqsjI0uVzC77kDDLK+w8
10aF+2ygLeV6su/2JgkbN0ACO0vvq5MFVt1xEGVwExKrdvzmFe3f243EBQAORBd5
Sfk0s/kj7YHdnToi3wnUQFwFS+TpWSqESDYaV0LVXRX/2DNJYFTZI30gzzCc80Z2
1ccH+bCbsMA6dkrm5oAjQhMhhRAP4uVJvVF0FTu4Ztl7C9TJT0z08clNiZnfDVgJ
3XbkPV1pLqV+r1n2IZ0wZj+NvH4OD6oaNeyyGZnCo/gD1AQbBi6JbKrhQ28vVnCJ
xMxl+2H7RL6bObOjx29xD1hOfYReHcDrnJDNeLRM5r24nYiobYY9saCOjvp29eaC
sfnaiMXV1QwkiftgnqYdoA/Uf7ZR/N2C3hDjFJhl7/blqL3GNn9XVOWIgrf9zssR
HwBV79Wu4jd811px6XbvKJDRwY48bx9wz7mNPabd6j1h0QsHt8LN7I0D7WhYl/CG
CTJM7osXpqKNPwfYZrHc301Du4FUTpyI7j8ee7eaWbYl/B/z3pnVpbTVLpGJ3ZXJ
fxGPROtRHBuJTFnNyoYi+1KCWqLNJXmkn7XmytUInGYTUKIY7bcvH0NjFdJ54sZu
Or3C5hAhk9/nmaRjS6pTLbb/b3v6UCDOO6Me4tJMqgeapOiWQPuUibMO0LAETyLp
xQLVM0qFjrMzgd0OIEVWgmu7pE6r6BkN6UMhrhHqaCI/O8mG6XcvzVonnOf1GK6a
CXD12/sLCZxjLn8PkgJWep2L0qxrAW1dzGFe7qO8Z6Dv33p9EnC6a0Wxc0Yvtrke
l1kwopnqB/4pmw+T8hiLDSS4QCQM6U5CCuOIqcAoPOqZWKH3v54mIZ741CPW7Dug
bfBnGzZNClyx8xrPvzIKU0PEjfMePFqZ9k3Q1YrwMFyg6bPW3AB0y17aF7dIt9qm
d3ZXIbZXnnSlc5B44oX0Bj4D4nC9ogjiipon+D5b8Hi/L7Vd8rUJJvfZzHIOlCju
2Z53ZDsgFhz4Mdeqw5tDxz5RBDCBePq1VsYpGP/Kl7TtXDH4xrohnSC9hCXl5IJ9
hRQKMGHL/whHqXCS3xXS1sbwT73exATDVrE05rHKwv49NS0hdVpaaBwT3YkyLNgY
tUEsVK7YL8pgdfuy6TzD3uFgvuAhJ9fKl+PSmXP8wgEklukvQrx7IUICBYuwRuUW
/BjrzrPpMN/ulm/gdCcMMMGVtnajavVue5gF7YDK+W4fnM5/IcVEiCakPNxskjKv
a+w/8fROHOQzI1SGjsKD64TuBSM5haCxVq+6O+WTiVxOWBbUxoaFAje/BcOlbgDZ
C+b5n5/J2/q1tEZjfjrOZK8GrUT+dEUW5b5j/1G5AwrWvKUwJAOkKIwqTfVdAyaT
L7gFKMf12CqYZt/hH/GeHzalnav95ZDvEYSLsx5ipaU8nosolZ8fdkEapuwWLQgH
Cx5jcFCMbhYW6gy6hxAMGGY19Hcet623CoAIUF/WOH+2lAKADbSjCfSwANi6ejDW
BNPAy3keFiWyxPJWkjShm6EY0TmudGN7cd+gRJHPrHULg2mb2B/EHKZS7JziZb60
oca6YCzg96mLpCs1M4t3+YeW7+IQct6AGdPn4jQhkATRDDjrbNMmaU73k5fBxNFb
PpT5lGM8vrZMf9gJ387/zVuNWf1d6zAjk3fazizyi/zuxB0DUSpVZCdNoCF8S99x
a8ZkNh2bqbsaJZbWSO9XailBlpWbQHshV464rv7zE3H20/nml3YhiXp/DAHeN5LX
h8/7/KnpMNUghzz9HKExS897pgRCpr05eXA1iWVb4G+f2Q93w0IyCoj2NVHBgCfq
8G9ghQ2pi8SlKmQYptc88QZtWr2OLDph3Wub2MtjtZH/MuOk8k9SGp120l6ito6k
gxcrW8LSbWg0zlzPMkdGaApDy8WXrkxynML0cnXSAEPWhv3FE2e4SmKXsm/xhCQJ
/2ein0BXyotlQ6GZO+irkOFgUsYhDvQW5lbk0t592MlKjh6aSpj7jA7iPjqgULG0
Sebuq+IHcQkYvb6bafIwmT91noWmiXcuP7h7th6a98MQOzsPOc2hSH3fr4ZuWDiC
ig56OnfDhwK5tAWo7ALXIgDB4tNChWidtosG7SMKfVKfANtA2qjfCX/03XQuUNjF
RwodqY7YesCOWMKvOw28MYzW1m0SVNM/7mVCy4b6gzWF2/u2cbOCwjwfNiQni4bP
vno+rYUIA2fW929rTVSFQaYjD3q7Co9m0qWitZQ1P1Onw+6xH65jYWe+0gQjPTZe
WQlsl2FkiK6WeNEMmfYBbWtfh8XlK2+oQ7wMzJJuri8nopxI301ky2WlL2b4Wpr/
t0m3R0N/UpIYpwTT7HwtoIbB1e0MupxVVhKrDSWvqQiBiAOzkrmEg+WZJLtXZVv1
zR0V9HF5WOXMrRcrFwH8vp0m9KYAx8ZcT7FJCpUqpqaM3xw1VStbsFZ7R/yGLTCv
puyiPwCEpf/8wiRUVbsJd8BJSkfVL9+68OJH3VOKzje4Ixp2h3ykOZKmKbCDxQfn
YiNei0RF8yB5zxwLzqjZEclCS1d9U1iJ2r92y9ft1Sl26H42AW5rkZf2y4adc0qY
yZv1GEDKd+/mPk6czMjGYfk1D1Ba0gy5TfzAKZXYEKbPbeXALN5/pH6RZ0rO8ixU
kk6U1FiL8stJjhqk8P7PUducSRjyaLWYkUjNnU6+lsGiaHfS7r0PC1l0or++aqUA
0BpFiQWPLpYIX4PHoG7xX+sQoRfUuCJQpSkpPhx939O0N70rzykMwwZDfY161ay7
GbbtQ0SEFBqd4PSuM23g7lO85Qf+QI20SXfMycVU/X4HImPFjfj2idg8sVijYjCS
b+cf5zK+P8uv6pUKAZW6D4nHNopOSzTqsf/I0dUCul55ldafaMjvKh8gm+76W5CT
7eh+QFt2ynQ5hez8haG8mTPB0iGQDWmzl1OaqnoWmdhFGqtYLVu97oAzwTBDFaT9
xqICOBwJLscdbeyCNdUq31+I4oJIac7Z6cWO/PtD6l9hPhbvE9l0xGqZhF7wxVj7
0P09C8m6/Pvzcd+Yr6hP6Hs6kAXN2TpHXVOsWk7/WDwSxfkmwwhR6TP7S0Yyd7c+
Syvh3aieINyEQqbHjqeKr2vfO89eD6fJU5GA9Evaz3e7fr1rIcVVHmKes9sbBSct
jldJj+F7O+o711jUEmV66SbzEn5XKoeNqw9McGJ0MZQxPj/vc2ZjYVJdtBovYd4Q
xh8DBojTdJot53Fc/iYXVJcE8MZNjWPh+zAtgQ0eqNl1CZipa2FAja++ioemMpq2
Qs3BNpq8HN0tng5zpENNEDXMeIjCJQIZ5ylMT/kePOGFrSX4itd3MmdK2kpD5YY2
VQWWOcBx9QIGMuaXSwJ/jMS2ZQS38CpPVi6MJq9hdXE7e74iLTKoMo8S6csepUfh
8Tt7AbLfkD5P/Cfd5G47+vpXY2OcZYi6yC60bh77+iIL7728MjdGCCCbv/7dHi9m
CCCjlVAok6GP0suC4RCWGEcBb3g8mzaOzCYJ93sfVVoUfAOLQpbUW0o76dAzjsC6
m6HFcOaK8fHnLaonZOU+n2+IlEMrKP4LlM59Xn61P5xmyTqdok9NqxYmwbovDGZp
NVfYWvI4pFkYmRCBOyRj74Rhf4Z/vTV5mmGwSLYK/zRAImw31cbIWCLPwrzx1+zp
GLB3FTpaBht+vq/EdYplXcPBF1bYMX4uABZpxhceKAdDQO1VjA9L3mon0Eh9JZKn
DMVeUMcilArkxU8SAp4r6LwODebpenDDaJNU+rKvBchdx0SB41/V+0XMEMIrc4Vi
vpGWZ8IM3wYQVcwijfczCRg0kNyStMvhF8/TgLGusgoZVJmk4Q+PeQpg62Rc2dlA
/MTCUuZPSIqQ+ded9In+NUHTBuepXYNfC+W3j1eJFiAEHTPeO/wtg2z+6Qf1djW5
N64LiL2yMo5i3SKUIwD0UrY/0dhTiekoy0KFdCekOdzxuQGgXEuR8ciOHq4fYxNv
s5mlWBhwK1VYY9br0SRNXDxJTLPge8UcLuM4Fzib23goGFMqUZaIhSVELdXttli8
+MP7tQ3g26ZoHCGELRB6PKLRvdxXwzTW/VAmGOzj1AzG6W5mrmhrCfUDGJ70pGiq
QoHv4R4qEibBmipIgeqTssPi223kOmq4/gl19nPusK5UhCz20659hDl9cXgKtlKU
Qdrr5fMgOLphAwRnhmq5eXOsMqiH9bb0bOzCGJfw1yoQzxqqjpUjIESdZdNXeJHp
EIIgCipA9/Sbo0F4n3tSyoF1PIfNcdpG2PjCt8jDqM/kdwKNVhL1LO1jSaiI+Hms
RTN5ZQ4vUCULe3ya/xP0qASp3zOpfeOtyI+4w33qfOKVP2meuS0SnRp0hrd2tbpw
rqjQprr2fY0wfgQYLLffY64ZIRrFffqRt/yqe4w9V2Btz96wHZAdXPsPjR+dDn+V
BMIzVd1hCUL8dnqzT4q5cVb9+uEP/ChyUVNdB6vuPvXV6Zl5Ofj9zgOnBa8wjc0D
A6156GIrziE/fcKPC5pMdHou8hS8ogC2xBzGcWgjiXb4Upwjvk1Wg1HbD+USO+Bw
KE7QBHXKMXnvQKTbGErplwBBVmvBiw0rChsHaB7Jd1cAeVf9EXQ5iih247P+UUpc
Xc76p16FTeBLZcLIP7lw5V9CKFfH7fWGifhWG9zSfAG9pKKWtv3zbj4zcw9duE5j
Gnt/RU9qhTw/gkx4fT3zc46+LlXPaZM9pGOBSWrLQgZMcEYbJ/u/bRYGScKMnQ7L
RTE++SxZ2b5uwnPUM6Gk7rP0Uy3jni0QAedZv+56IJEzT003NWffKUWYQ8PXl2MV
ucHNx4OBVk3TWJqfyECDdspqSivkum2S/uw49gUxUlaoLUKvd+QWn6XSpGZs2rze
3UyF3etTVUZNQtJ1fZWRwrQ6bgT3Ryrn1kiqrh9H+Dxi4xPyfLNfzykc57YB48Hr
5MKqUi1UaJT0sQZV5deX8Qx/354e+E50z4pEaXIri1G3+yUb2iqsPlYCLhNBM+EF
68hkgkDq8oxKGHKxZt0eOtE/v6gieSV2E35J09fStL3mejxUMowcaNYfT0xcIdS6
MU5isYfL8idFp3aslNCjxBeKkeNsjo7S36lp5vhTGWSdOsLZMgr5caAoKYJLvZS8
Q9CmvX2OJkKUfbCscRr7bkg+Grlr5/X0X8g0cqFqsomP9AnO8y/ojJY+8jcvH/E0
kKpSG69V9jEvlv99RF2C89lrjVXo6yLSp8JynN/7ACqvBZlrgyv1M1o0HznPmaKc
+x9Yau99C+/zrK+NnNqL1rhgOeZrB5x6qbXdsjnr1v3RLVWqROYQRmkzXIADq/Sl
tSM1P490tcSMgNkheHRSWhKlDGyP2tNJ1CgwAzNfd5X017KG9oEeRn6pVCFSm5Nq
l63hn+57f2sYSN+wu34tm7QhxFORw8WvFDyZMTiHugw2YP2wNFv4c0F+tp3v33OQ
ikU8zqip9V72oQy4c3CWWhfELh2Flp8f3XxgHg+Sya//3LmMLS9DPc0f1RJpyzT+
xmA2ukgiCEc00yTCaZ80Ya7LlGZA4HEl21/TodPTEKbuE4gZK82Wz7+SzTxhkGKE
X180YP5as/Fe/nx3Tc68gZp7uq6sj7FKgS+oHtfLVgSAt7DZnhB9f/a2/OjoGru1
3XlSlgyKdTRQ6dfSrxTQcjFpF2Wa7hawohkB11CRN2NJhc3c7TzWSbPGj7SrHZPU
OUwZlR3YjeOc46YlIfkjH3WyzH8LU9vOBQTDWeSvmlrk6EFPZ7M0prMfwZFhUHea
3l3JnDQe+8eZ+NJvivcnZlI2tQWKSkSBWt0N6q/LhClZdEL7YqXRADaGdscWEL99
3l+bjK2u/xX84O2Q2cBLK9SRstSDzFDTl5EryhJGJS6t5jetF75HmTLlYODID2yw
PFfn2Y63QSMIWYbzfCtvwWvmE2tRgV4bI1Gf65Bs7Vc/n6zBeZ3BnrEHngW9fv33
3YsNsdqFQmdPbrfsJTeQ8SabBB7LX6l0DGo5glmWzgrvF8HfvFzbkRHTLkLbL7b8
24udJpaHgUL3+1cdBc7OpauTlFkU87uXWXqRGmeSbxqqfUphp8/KC+mjmYgfETkQ
ZheOkkZpiZt3cwZbfC1nTiIodIPYCHKYr97riKhmw4gK6n5l8cxdh+QAY8wPtILx
RiyHwfUW8N1zSAyNnBQvVGsGaGJXxBFxpwmnZ/imkawqYbOQwUgWErO43mp27Ewb
9eD9G1B9jUO6rR6Upzgps9A/fwOCDoyxrVDdndRGWWUbaVwiwA8XQ7s4h0RRKfIR
B/o3M9oTYr8dw0fPGoaxSq2ZO05wZqpXXFGSujLg/a6rcVbq9OQDGInuKDD4lD0C
8tqqsYQz/dpT5/9fJwN8vhH0c4R6A/jvRfMu+0tYf3KINIMBbgq9L04SAQ/xXklM
dxu9wxddajJHX+Y4DRSHKGWvSa5kloP8aakFZ6Dl0Fi9K7oW7lWaKFeDYiotTb43
r05PFUjFWZvSoAO3QSoAaotm9fqQNjEcg+HIyy+zr7elmZqWpbuDw0Yhw4WOPt1X
B/SZ9azB2wZYdtVk2gp1WUUflGa26t1mVKQv/jLItZtVpL5kOaT25k57MGAxp7/r
dXwPhK0+cuAtioZSraH/GcOmsXzBjK91T/jAMPjeWTR7J/jUBcmVKelmq9v3Vys0
sLtMTPVypzkZ1qb0G/03gavmAvClyjaKPUBm37zlDoAhNU3wflIDxcL64fQ4Yi4S
WMZQjZ+rW+iNDS0twiR2ACwkQb0O87KbPnw33n84uBOY0ooe8qcnUy/Fh1yV+Sdm
UwCSMQTFOUy1i4c3oalD+3VyBlsPY5dWoVlfBuUk4/ynfQG5rjFhzbU0RnbVFEWh
2VEc/7eXiH1Nu0+ucVDFekr70qpwaDqgES7hQNclAkOwsJy41wqlkPcReoO0FGnT
9IkUb6PXN9HZBCbiRXAOF4zxnUbqQVKlEPc/nuFI8oncQ/46yds7wCJq3ZNKu/uT
m0qxxGn3sf/yR7uIj3uUz/TgHo94MtNQ0l0RaJO4SpYdx+c7MkuBdjPEurBePGk3
3xuFt3e45lOYbS9abha3m1ArGMgq0IfSnQIohVwXFOK+z9Ho9kE4hf4OSzo6AwoJ
a9f+B9hq00sq/VyA9T9lNREFuMQjLVKascgidiyC+D69KIKcrNhRGo3oDVJlFIUw
1gEfm4F1FRX+tCw0ECuSz7x701oeKKEENBVjiumFle4u7Ux9VtYhm00Qp665tAto
h5GvVeceHyVvzxUyg3SV1uQT3yfL5E5zYRU/S5ES84HIlxkwBqi+B7RyKT4t9vcC
h0y6Jg7M/KSxJ58zgyqKOlWwRoKzDeVCIStqk/5rb0tySfCWJ2B2tXjnqXWyogH3
GGU5e/eiD1G2KtLIC4DZSVqs1OkZncX0CKm2RnthpgSNmRQpdRMAcmySqdUjahxy
9dyDt/SmlM3Wcn6PEue9pI/YkBbIkjl1wAPX8W7oM2ta75x84aD6GedMM4SsUHoM
iK0gCbQNbw8wndTB4sRZo94WplQiibcHY3ngi+mHJ8Aa8BsDsHp2kgUaKpMWQWp/
tljMrchgPSdI8cpaM3GLG9jOJm6YQd1o4QREFnylN6lcomzyYg7wpzxF8WaOkdsh
3XJRhTnl+WBx7iq0JdgsV9gwHzZXXu/G5pTAGJBTHJ5MJvU+6I/4S9isQRd0GDs3
rS4hbIP9iBqOM/5czPZOJtusatmGo+7YaBt24BO1b1OZ3YUii53z4W/zk29TwwaO
yv0+015fvY05kxW8zwR/a5LNwgNMOPFbn8O7PyGb8vkq3r1/a7+VMOHaKt4/nD9m
FjSs3avNjqU6Uruo+1f2oh/Vn8yAxNi/wTlHbMnNDhAfwt5HpwnUXujJtLc2BxqZ
iWBY+BrlV4zA5ocj2ziczqpRmlsWKx2uWCFMi6jMhviSTMpc5njOmjkyp+ryU7Pm
gP+BRps89mdAexLkKDrTF3nvQmeDEG0MUgEYDWCkWgs9xk2T4sO+aHuH5lYOVzzt
kKGY1i3fpYWzBLiaVMyPImaIOWh3AG6ZlAbCD28Aj6PN7gUWRxhvxLvRPgKVtDAW
NIcwhIATW85p5PxRfgUdPYItzxuAT+iiUPu+zNYjBdL9MYgWW1aOeuLCQOSYbBkw
H6OkqNx/Bz/rpyeLD7v28MF9Qb0OoazFDnK4t58IP0pKQ8xYtjbIaaJ0P1dvcTuo
2IHweyE1LT5GkJfB7Eqdx5V2FO6oxxwnZEIkYCsRIetYdH3lZnaJj/WUOEN4fqJu
sFcxOyHcYyiCLnKo0qgJ1YINMgz9bV5Dl3dgqhWsmUScuuwol/LyfFTeC3TvacE/
0ikqy28G0PS6ym40+ADkob1qj7wUdH2jwPv1jKuCAJaIzdglBunaZnOPSgvWnn0p
LOQRiHQWeZx3fEs/Lmez2q8JX4ak82rSRQzrY4Pd1fSrst561EG4XV4oIFCrd3Cu
K3L3y/rTvjcnK22LcUCv5XBygGKpOc1zyXRDvvIgGHdNF9iEwPk/8iltW8+xJEiU
aJRSS9HBjpGQv2tizegx3kjllw7TeXRGitkT5DEWVez1Fgc1bjVh91PmHUutkyx1
yAOTBnJjRjyRhxdGX0q4m1iCmCF6n2/fHRNuj/oFY+NP3AEWcQJIQgZDusrp/R9M
QkE7ATSWHZk4UIyd8vR/lKqO8/+hUCHLx+cem8I+5jXHiz8fT9fkImeQmxu65plE
WGN+ccqpRjUpNsyA4LtyeGunusMZbxh75DVjUC3rTSHL686TV1anMUeMC01g2qup
SaW2Js7K2L79yrX2eMDK+ckVh7q/LPMGp8pV3YWnhZF/+9nNAnXjjyY6eGZ6mf8h
N5ffuIQjR9sVPWikjAasmRe7egas8HvQga/1n8qM78wWJqRVt7JDaKTHkxX3DYjD
V9U0kFfNe2a0QscjTXtziijHmWWV4loQReLezkpWUMlsPngzorv7FbZy5sBV0meG
+HSxyI/6GVL6sdmZQuIoxdJiScT9LKl73SJss/RVCz5O5DhZo9TuNhqjyWph5VGP
xKKOa9U7xAxPq7nD3HWFiWlFbTDusgeUcP5Dcp9g+UnZdt49AoSQo7mMhQc/ILPr
4J41sekYAeSvP/vSTNlt+P8kEL6V2xx22CoThv95oncV5OL1NxZkjQMhd7Z/mqv0
l0nOjBgz+ZNnza2qmwUKxlUD3TXyA7aY2corZ2OHyD8xN6MUG2967aNC2YhZQoue
u1PYUAhZf3v/d9IbMaB9vMv6tzv2oT2SyJS640rV5NM8ySN6pyq8/02jf3w++uhh
n2BX/P+3y/ouk5pIVOskM7kHFNZBn/abH9q9FfMJC29MG0g5wsLtxpLEMwl8TTtq
vse4AG2hc5gUsyVf4cazE84PMM1TjpWwicaAaeiOTYQ0p22rupa2Gq0vx+neRiue
nq5YcjksyUx0DS9mZntOtGEc2pOoB6WAp9sOI8ZW8nyHMMOLaspAZCi8YZ5POmxE
8osOsHbHuhQqZYXDB7Ydeh+thQfWQ+ZgZUsuQAql/XgsVZ7l3BOSbLam/VqZuWR+
tVrsQwaXh9Vcpy01wn6MdyGH1SqcMdcHdToPj6lPRkm2NH4+rE8PMXADLzp+wz2c
Zs1zeXrloZRcDOJBIBVUvQ0XnZ8FGtF+UhPUCWG2sUIdrMqaZPlxwyjB8KGKheMz
JIOvH3Zk0v6vkWYiNNIiBrh+aPRvIIywcrbfpGH+NvFb/3Tzunn7fBs4l8OY+juS
y79gighMnO+jaPAoZD706jQ1EsCtZtHha9yWY3K87qvXwXU821Kiw+iE0LsEDV4C
g/MJOk+Um3qNmZMGGD6gJSdF5Oalj/FS5aZrQ1siLQ1rUsQ5/eAji13QTRBLj6+X
Y4D0Q2JN2EVVn3bU/B1U6slCf3rnegu7d7SMmrp7TG//zfwbD77nbUncTfSXO+Oy
poeBGo72x4TDfuJdHC60r2gggu7l3apimk5FQUBc6MHAEK+KGC8/g1nXqhaNtwdI
rtBMPku1RmXIqnaeWrPFfxYgfTNqXNa+yNqMCSGJqgl/58lTGa2UEemOLveZImXY
0g0ct5Gm49cxOxU0geWUzMwzj6hYWL2RmBvPcluqTRgA0m3NCxFxGAfZjmeQXSnr
X97yLeDD0m6WKEAz7tmASpZOOAiDDudJoGA0B2WEdW1GvfOIZqZSHXs4q8RIoRi2
HCnoZm0Kl69lvoaBJvZ322NbjNBc+FP7ywRmDeBdDSJRkJLf74/gKUymXFA9T7rO
/IbY/ayUg1BWtRJ0nMxu7dZDuwwx3HikoJbEZ8XO9DivCOEBw7RcW0HEz3Y3mX62
FU9ojGKEh7Ua7u2X+AMZuoVJIsdGgR4811mMbrxYlDKWTZDHZSjE6REX1ghQdEwm
t2PmWpHwdrwpVltlj/QVOgJ6UIISNy/ehdK28lan/V/wxqEIZo+dhB2WBFw7XjWu
R4jQBsFY1iytaQpz+eH53f1HbI+4aiiM79C6iaVv0WbVNtNSxeix850UaacyqrR9
cU7cKzUu8Sspp4ezRDhJT5N+s7FOGW9QEzTgx5SvQU4QBg10Ce0DkaULtRM2xaZQ
vYmQirFonsLCqp7ORxJN1BDu5zr2PbbnuN3lX0YAhJmfXiTt8vnX4n1z0g42Z/O6
RDoVNpOWq9DbDX6fFerKD0KKIOFUjjW6SUD3hP2v3VMrOlIusaUbQF5iE3czQMsz
A8ZYBM+QowYjAA9EtVlJkfdsky52qYgOFzBJMcz4F+2iHEHtVz24Jmc1bWm9TToL
V3qVScc39NhbILQh/981p8LNBalHGtBMkKVExdRR3Z9IyO0enJz67h6NIaCFfURQ
PH+yx7xmQsHHGbjaGwcG2wefRFAdPvwpX2zYhuXGttZ6ufxaxT+Afg3sGrDvIzUE
it38cAvoSvyQoR1obhXHqPSdsae0+OSwhtOBnTJRMUCMLgYtCbHCaVUxaCHqkSVu
FfydUZ8F8UCWT0WxbheYhS1oJkCHEKSqdM+719fvIGdmcYGIBDzSuTYmxy60iQXg
WnFeHvYEb8p5YuecIXmkvAdkwlZh+Q6I0lWniVJENcuy2FngkOaJ2f/oWSUhK35O
JCOPhyS+oheeV0qaxxk8FeWWu+EPpOaF6Q32TjhUNm9jgjJpTWcWXGF5PIHgEaxX
5yZ7KRXj1QGg946g4vQO4JtxvYgfs7DAuFX9NrEG3dGlcCLHIHZTxzZEDhAzLOmt
yM+cdz+wfCP3gnctx1dH/WnsMzGJAd1p7kMgejGlm1GB/OMJgIneE+RIakuufZfG
G3BEHN9s9hsuQ5QSuubXfbGY4nNL2Quz4nBnIBL7OAnbZpYQuF+3VGKWjuGZREui
4EzbBSleM5PmMvyixCdt155kdqmXVWs+DbyrXGswqaaAhfIcCECBJZWScqwwRBuH
T++PJXDAUF1occ/qXIGgtz5DnbZY+2BsxgswebRc0xgw+OmbDsSEqYsbXlo2RlS6
mcxn/uOdx+3t+rAXYi2LXCq0A45knTIvtaKPCYft4MLNO4srdx3P60H3Qt287Cgi
ELcl1KONy+eDe/ejJAUs6ASSgnZSy2uVWnxdVuNhRsQB7qfusz4WBUWukALNtjHT
e8fNPcEzlsGM7UzySdbdKh5R8plDxkVP24Y6hBzl7R3KxWUyg6p8aUXSD0oN1C0z
haJyoeFkiqs5gxtae4yih/1WeG//Su9JIPIVP15LM8m4NS1wxB7lxas9ayqDSbnm
V345JwuH/ZvpSE32R712Kc3A6ZJ/6hOaOR3S1V386Ez6jM05NPjWlhkdHci32yxz
Gs+CE/WtTtY2JW+77taRj8WFeYbPCtYMIGEzB1uaQOVTbR6JBRULEbl40HoyA/8R
zqrtTQ/9hlazXobdAnyM1RTLxOVjjBICJSi8aZIiBwioAVmI+0LFOaW8a5ztK+C/
N6Z6fXK44Vmtl17i9NsS5+hsUzo9aotDYrB+1RUBlkTlH6CWy2jV6dhpG9cyfjal
to8yrAa9xado+LD7kT5GJ+q2UW9cFC5085/7WVWgumWFFRRYKAJ37mH9Ti2fyAIR
/i18fVR3o+TXLahjjDd1hiS3q+csEqItTXnpyjKJh+LAo9ZgmAAYIT/+ti9Yjbup
ylbBYa9LkuHVcoYKtP5rGjTFeZqOvATpAlY+MObCFjxu9W4GglHG603EwNd0FkTB
5M1EskiVL7I3/jnC0E5aRtdS3OXNjoS79PJQgzM6C8eL8nkA8ICtwXgwbM1VqU+B
/jF2L+mSTyu5Lztap1NWZ37npblGeVStLxQC0QUML1gB26XUmHpYu0SQJLu1Fe+Q
QD2H/eJE0qoBqHCcDYLaKwhyCOR6eJW+iuOshB8Drd5ryoCJv/NM2ItBqj6HbbOE
TUKE2YZB2tdIkxRxi/6ySP2a/rFremMA8B1lmnA/dm4bSyhEeXE5ZhoW8GvsuMw1
tAtQ6B3zNcs+f++u88+zdCHkrAH0COIomB60vY45sN0A3iVbofeIy4W3reDmr9fS
t/dM8ZO4uIqomgZfoe60r3x5mxDS/18G46JKcE2AYKZzqy0omSTUsUpSI7cWfM0o
LlkAJ8w7r2Xp3QWSgUn7bz6rZvnpx0hf9yCYuBC3ZfdPtX5F1aDKM1AQTiE7VK1+
UXIhXDZ2i+Rftbs9ZL9XEKSWc6VmyWKwt4m5uvHKhbPeo6wXXYDHhEXbltbwlKSk
wzWRvAm7YKZqQwlbi+P+sYI+PtR+q7tb+bRwh+7hh3xL1ew5M585Tn6aZ70Tv7sF
K+Po2EL5iPpi2ZBq3nNTUGr0Rmj0KYeWf8cw7PjM7TvCdiFAQolbWOooKuL5gJUC
8gkacUVKyOgmAm/E5D8JYYTySklUs974+6rRLFNOcLFQKqXC/PACqzoG2oPVRpUq
bRJkSAi2esRNogNjcCODYFTfc8qSS9yNarcRuYjd5/lZic32jgFDwQGGfjgdYfxp
prUW6TMkfRJ2xLWGEokwgvUwGDddR5f5lciNv476Jj1UR0sApJBHAYiHHdff3xXx
3JMDdoy1p1JKiIOWwsU/VquVDmAiR0AqH/4iVRfMX6Uzng8fFFOCLM6o0pksgMo5
WbhTpl1q/zEOLN5eIyJ6qVQhzTJpICYtmFMNEVkPLAmc1yRbK13ZiYwGpgO9ls9a
XmGdPja6BFnpob6dYvFWv4ZvUoyAx5Q9D0IlpwO97cieTBlm3lD/9FLypEvn5HyP
4E2dIvjtMNxNQGvXW8fiL4KqiByksNyRkdWzRuB7Awk2PRdvuy1ZoejNfUUBPNpl
FINhjuIRwDlAzUww9v9MG3MdZFlxEzc8zveabNf8lOlFufybPdi8nk4NceG7gd2j
DnRIt7KYTBgkjgC1aGC3qrvJ0+N7tjGZ5m20ECmvLzLxfu05Lo1gmRwngpR3bw+R
XMI5iNZksKw9cneD18P60Yal4Lwut3Hw4EUn9UG2p8oLdMWwzUum/8WvedYu33SZ
98BHG6gVTHSlhfbRS9lptIw6+LiphMF5G8PDrUB05O4LE3bURYTo6+w6xrbhM4iG
k81A0drfh5loRnzHhfhZzaukX5+WPeVf/SmPgIRpt9fOI0BDAdsSlyaLyBDK7fLv
mOp/L3fXxPVp1+Z54veHLdFqIWWvVPLu6Ydpmw4fuohYKQPO7DqL8uZGw+lymZds
oA8QcS0SNSFVqBu2t0GD04N4bDyZDkg4rgQvfhWUBmZQP4FR8hrPkYF5TxY3T2Rv
he8hytQh9kcIDRZiSaN15XSTl/oc1V8/MEtUt8F68FT5wo6l7FlFkY5paVULevrf
vp9lD+w0tGn+J8MluXXLiA89izZ8VNwzhl+mzH4AUrdFTE6pWmkQFJz65r71vpAK
OPDRctopqDRzS5sZCQFnWGs/xnk+WrS5tSAPf+8xwX0/NS7VB9H9fSo0ryb38Nt9
P5JnhF9UND2iNNUgY5DNLbmIL7GmbRizq8O1d9SMyKxrzHXixg7nvPJbn5QM3hiY
ukwLhlynNEe4U3BG05iR0uwIV6iYPMMmgEGcOUwqxmWpXLy2BqpnenedBIfYNkiY
zWswSsJMaLnNHiQWNMiJGBcUAQ+Pw9ZCKChYuEvBjPEKfqdVF853DhztkJt7mErU
+UCETMntv1GMf2AXoFO7+nKgfjwrpR/rCOWj6ADPJjLDv5NleezpbgS8IY49KiPy
IjfKvPHYNQ6mOhyPUhsbjUR+lcjD0on9g0+esjlLqVrFxIMbYH9T19nVPx5brnPm
GNtfgxhbDLZ6/NIlJJcUM6PW+OXXBWs6QCe+dfk7JSLj2QtluVPF6WgbpUGhDUIK
/c7FSUOey2BffNYBy0nOeaKmpl0Fd6DQfYjdREi3eQ6sV+lS41U+sFTRTVEP2xcJ
2F7WBByuJkvjWIBtK37+05IIcsrEX3hvQTLHeoTS3aqHzwaOFZuXn2YcPvUy4NyS
yWd6ItGV9Rz2NHR6zdDGrZoh+O8PGNxRXgot5ZyB7IuPUb7ZvqBU2u1a1coI52qC
xPwqd1rvgSJwbVGf/Qq54kQ8uxObKNqi3fOX81hqq8nhwnY2ILGiv5JbUHhVbsSW
A1rarKXbcek3mlu1sadMeBwtV+6cM6EfqeGKS2jYgXp4zdKxXT5xbi+KhhNc/atN
BtK1w3wHauqzZMIrls2A1C3xu4bChCbo9W5ovKjmh3avLDuEaYxueKKcT8qSypXJ
MfKd0+lpK4C4O60jSA6H1GIT6qDXQ7eDe8rb6lSKLgsz42/iu1Edt7jPB8gfBkoS
qv+mDEyllZ+jbDINonQ4QGsj9FqDIWfYuF7Mqa9S3IUX4A8juFuhjPV1o+vCpXMx
by1XMKcoMXpNOCxMjD9aIz16hZOoQ0gKZn2VJCoPMXJrQ36klA9H1wZWL2A7og89
UtLyEXrN/2py63iMGIUs9rqyug/U87Mv166SVSEloaSv19KUjm/tT6YdoBdI7XkM
/b2RiJy2nE2vsvTROJAlaALZ5HaoMzl4O5IFG9uN55OBFoJh1tozS7ELiMpJlAR5
sDNW0Mzy2edyN9F+mQtraRaDVFk3ax437qe0AhPVguQcp+ZrriXnBbQiTwCHhT9s
T31iKZxnr3DSE9LkQLZIzLgZthgkLcD/ED+DZxDCfhlYCJnoQD/8PS8+cmgMLT+z
ke8982auC+CxLCpE48W7B2zuW1YI115ah0YaG63M+eUPRlLC9Geclkv2RHFQgwBK
gAXnWIeknK7W83A0bJmYCSEuVOHbhZsbc5kNF80BSxZK21gSn5udvvaqBOyg6Mwx
up0JQFXdKEV1sASQ40OvPD2d0y5qlajLCXeV+0riyDrul5/9nnp5ZrBO2iM8hl9C
fpLiVmJj7aN6LpDbinu4qaPnphJz/tJdl7tX1hS7mD5LkBD1tkoJSDd0+TctkzQx
jQlLwdSTslLPuvVcTmSW0BtIcyUVolEHn1B9Io6cBaqzM5Wbhu8QKEY8VCttahv8
nZhAddeiRydqDBDdaLoEuzvDBRjzG2Rh4dlWkv0jaiKhmEqV8pr1q6Q6CqNsSv55
6KCPyFrcVOlXmMkrgg1bEBpA/zFbE2zFW4xYc+dhQ28LvXlCAEw9sH/pyPPDSnft
r2xsJGON2HksObISN6xcp9AoBqVGMleZsoLjNrvxdpMg8bGlL/G3v2qDayX5pRW8
sMolnJwoKlpAqy4TeiXjPPJA/kLALSysUD37/WxHAMHqfL7XSj9ORtl0igTcwyT0
MzkU4suz2XOAsq/CGyXVO6RMflN0RM6aKneNEPBqMO6qmmHekbJwPrlSY8C8QXAI
jHrwyzYr6CIJVcGxvx3CqZCZyuAwPhLIDQQkJrYeRonB+FMhVvJznkZPv/3gHP4D
WtOaDHOsPZSrKF7+NUJPM5DSzLY/nYlQBwOlzZpic8FEmkg051Sf7KBQN4Pao4k0
0yhnl7MK8zSNM5It9iptkAjFuo/IPUXWPDxie7xb8VciGVDv43k/BgAZ7YE+FT32
kwubvud3jXevU6Q76SpNWVcStDzrsVXZKMwlHi/xDTjdx0yko8PiQuEUBgQY2wWI
cJxffAdTJK4QTs5I79RM2L6g53GpusP7Si6/dbM9RRsWm9xcOSJENCzfdDhluh6v
BinQHMUYp21UEN0rglqvklUoIpNTotR5Y3j1+9blmFwEWeG5qEoSP0hvJsBl9iST
Rp9HlW/HUiN7Zgu+xYno61ye37grswWcsTNDWpXBbBJWxzKKwKU+g6mrHliAT/3e
35gRVpwRhha0PD64SvoHJvS/1p9FDUR5tiEae/cgzBakLUmUrDZ6lroVCGENqgY5
xwxOWXYcNljgntaO7zlAnZ0bMwNiU+kH7OTvkDkBrObY3S/vX74jQ8b5vPe8VObe
PI1o2CYsxwoec8BlgqDweqCPU60O/HYKpOv4abBy38tkhKmLa4DKjCZ0QQLptdgN
p9mlx0O/kPhME3eR4R1RdaNzYbBLlqp1BspIxP/1CVtxgM+5Bsn7cn3HNVvH2SAU
ducswAWgSwM4N3m4DaUZwDyplD17EA3Lt6kJ1C0KY6AuAMZtipQfL86B4EB9VPbP
mWLaNOiNL7hhG72xpCaI2SVbnm9uFqCQ495VgiKEyAZaH/pA+NbivIHWLhoq3mru
hJqrkjwTFJoGYQsNAfx7ZCmLiC9BEQqyv1p361bFpknPfCQ67X5FgIG1YCKI5Npb
auJQSbPWpx+NsuDChdWYPV7W8JVuq8QXm4qFqTCo5GPBKe4dOvfNc7bNKtUaBvK8
3b5Issp9BboRkhjgINYx+HFwIDcX7HnNpvaApPBb7tMm5wRAsiWK2THm8N3GnO3i
/TCFojSqSwhOlHt4KURAAmEM0JiDIDwhu80vG/EcdVr9uUY5MeX0MVHuBnC6hFRk
e/2a4JQdpPOWvIamDRjjqzD6TKB2EVOs03lSzcu3OM+wsjMzuFUtwfi+VmwDgiDa
J8W1OXy+uR302s3cUphwAr+CV5YaWFylncoZ6AQpKEMLo9ZUy3heVLJAIyKQ+FqU
ONwTw9to0sPc/ViDWcZzrZTuQGrub4W9/EEkQwS3hkAKChdyLLA1C+Qnw1kkznWt
7R3IUrja2ziPZelRT4kodoW5ND2uJR8ctM4H0rQgl/k8cSWfD+W2S6UPuUoit315
dcB63Mg7H5/1UeuWReMWOWx84kZdZqcSPvW9HUPWoc+TQBUP6a1trR8HDYm5NlAl
7+4ZaR/YiSbPt0Csm3I6T1PC9VAXieQTSMS/8Fk1Cjw1JbYEwrBmGxMtZBzerHOT
vemVoludPWvUQnBtJZyKXdxqS3jfmL+AuaKYVSW+7zDUeR5jtpypx7x92epkYTwq
Rx9b05lhAc0tsZCN3eyxbF/rjSKkrA4xSYpCLBt85uFqq9OziPEYD3UZlcFbztjs
1myK0nnSHw8yPKbVd7YDpn8k1nWPR9y+EZ8WRzNcNSUaVTh/DdFetPvYCB2nSzvq
MbxJPyLc+n4SYWqzgOSskFnsbSgm9kGLd8Kt86T1m8ascaD79phjJ+yNI7wUtUqm
VjfZGqNHow3CA0kxE6MmU38zni6M6QDtua9Uf2T51y2cZiXVTFMb9TG0mEg1VvhJ
XKOEi73fCQAIAluw7SN12ILuKXIgbHY50GcfsqpFtija0j9V9TLrXqfv/kYI3BoN
Rh2XXCusV+snR/SKYD++/8zMyaFLRR1FNRC4RI4LZ2fmMg+EJ8BRrGHktEyjWE/8
ff8BS7xWIHdgAkU4tEbNo0a2nLRO5ALDI3OUCQfuqXGWU6ZRuBcJYK6rh3lEdnAD
YtT6KYZSEyIXwwkJVltRanm2q9i5pd9w6wO/agzAOwpssjXBoT4q9O+/7xCe0JA1
P+bIFyrNp+lHmST7M9vTWyu17sP5Bw0Oy8jVKZFX7E3QcsnolBUySIR+kO/mwSNg
0LDtyZhT8m8pwBHr3Fr88Akrb8DtdbQG80Sz4+tDgv8ySxusqvwXmOoiBBgvI659
Ada2i4G+dAZg55l2BfDX0cnDzPRacwG7dKJK+lWkbELueiI0IaS0wIuNnZbqYUee
L1o5bS/9VotK7yfYVzPsQLFEWy1YQqGaCgK3ZHpyIe/GhZGyqMimhBCPG5FOcjc9
QJewSAlDCD26x/AyQZvWj67/tXM6OIa3fzz71pdoJg7y+S6AQdia+dUzcDgdb/re
mtBnhkB9dZzO+aheyWaeWT/LagSdKl9KVMOAgKTAFVvPZPf1JyG5gFJH/01uuq/o
yNYJTn/1E1msowybGd+iAW36QgabqOPqr46TiTXbiR9XceAQFxNp79JE/hynXKKK
XmqFdrtTQYY53P6tTOjW1MY/N8hpSblqQ79KPuj6/7JfhxMcCR+mh5+wrAkMP57q
h8oNTPTxeYpFcuyXmdcBvI3Uoye7a3nC7/O93tbwltRtKbmnEClC/+/xW4z/y3Cz
xqcJSk+CYQsFIYtVrjERdAHgVyRN5w31q4gU7xqzH8dtw2QCHDqHyVPwXGqksILS
p6G+hipludZij5y2W5VYhZQbEIF4IGnAQPONEHXAQantanfjBEE0Y8mH52HY04tp
SMb5Z/d29EriXz/qvbm0977zHPvk9W3s3CopBWPn7YP3kFoxwB3umnnvuLNbU46F
73YiHl22FGFpRHMbL4w7el6wSsL1y3yJ7sKEt8+deEGJluT+IjHx6nUpvTySg4c9
qXZ4yATCcqbL729H8Hu+ffAEGmFTxAfTCLJ4ksmm8pOj2wQiNR6sG8Aul/6/ruHc
8SvUA862JMrXMfAYy0XcTL71lxZXfhj3JfhnKpmnDt798w/mtFDnd2OrFgnwNjcf
LVJJrfr3XKFUla1sa/oxsUcrzGVVAAl4ohMuDfv77Cp2xOxWj8/AM8RzDIB3h/Ga
jHlgmzPVNJCIQut7RN2ija55fZD6ECU1ruQc6PnRML1dROJM8p1WLkdKz6USzpG/
NPbLJkbaJtbF3YMNOwKzyzqGjGsAjvn+QnA6WxwOPcweRrB7o0oQ6me7dHJHSpCK
SbOEvDwkx+jz75n3KIKTGcDb6s9TubcQTA2Q/n7IibJtYOTGtB3/c2u9khbNwRES
H6I3tqVsDY7UYu5saddjeCZMXoqlKEWKW9JZhsNhXuWnFJ5jzW3F3Id66jHvg+lW
ZesQFvOq8PFbKNS2v3Cwg7eoDVvML+4eW5NU1JC/l3YIHXijMBzX7Bvyaom5rO08
YSfCTgYfOBLrdl+rSyOFmTZ8XFABLGySDQJTGx6lnpFYN3QGCEutiZ3EP25oIXW6
QGp9lg+iCRL5FCn6T41zASFHc+usjoj685S1QpuYuK164ZmAkBWYYnNdRTZGGrkq
D1T1BqtT/OoXoIqh/wwWHKBBPTDUx9M3/FY8JYmejFCyqhP1lG79qMPvKeKnIPh0
V+bslNLA0twUE6D99anX5079BEFXdTwmVD1XSOMrbfyAbHJ/JDZGOt+76p/9T+L7
eUkjSWCmGY8kkzA+Se52CabPaohBdXgAhQhB8IB25+gfdoCeSZHy1pF6jCGUdLvZ
jkzJNYNlG4muyFaswL3WRVOu5NMQmdiq21LNI80NZrQBqe3g2hexnTBJEYGfCuQj
KKhuZX4FwqKC0QMqVJrpuWT94dioPwMiFT3HuB6xrv8sv+K7MLKnByByEmSTWapH
pnFmGtXTH3vdrPaexX9Dv3BdjkdESBJDnnuM+UteK0wB1re2je5ua3/AKAXJoVdL
G0rT/munsLQj+A8p/d8KGQ2Gb2F+Vp5ob9KB/hUjWJ7DXMRKcY0RzWoh3Xdofj9D
Qj96RBg1c109QI0PIZq2BmXP0EnoWccEzi1k35He5doK9Ju/LGgtOTJlmaAgc4Qr
tuDoB6zoOJRwiqUt2Z+LtVSGogHq+3EAwVJibFcNce9j806fU2SFXb4tA3foBsnT
lIbWRnMNeCJBGSRSt+JcUsUpkhX6MMzBzDxqh6CDdkpvapvE8vJTAY1W/uJeUilf
W130XSVxW+uFceUFoJKmVm9vcfiH07H/s++kxKJb8ea1GavcrNIx+Vrsxl8bqCPw
CykEdwus40CDOf/N7z5oRtsIRhXKuWAabWF0izDOO/6+y2IEsXY+L2avWzCVW0Gf
PN30ZsvP0PIMEl9SI3itIkcT3JAOsmb95N0WUz2Cd3NU8ES1rfibCsWjpbgHRzjr
XWkj3qdPcBJIWq5PUCbm45G1VUhbhCa415W1TWd6Bi8IyDQ0Fl+rYIpH0f+sxcrm
CkLf7Az63eFhr5Px0Q2l8Fiyj7ekbtxRDr7mJ3ovNnvLztvi+zdlKsOUZ8EtjFbo
QJVNxOTSw+8geHkQqiGuLWipV7BQoQu7ag2r+lHd49RVYZqCCKVvg9bEday2hHfz
UR58E5q0MzBHxsW4sXaZRRhF7ZxVbcx9rGe3+3H1nHHf9zIi4V1M0K64StqHK9s5
+nZQnbQE4nxsiIZLU6waF/Irs2yIkOsKR732V2X0iO8cmgzHd1WecG+6a69yZeQX
E2TOFJWpMN4bOxS1zsjQA0JGsN6fzRd/nmjX5MhBvUbXih+lbL9+6LuE9rAIGPjy
p9bAxm1PKUPFVR9G5RrjE5O0AHXYaZL891PAPy2nYJdhxetaZ4oJrScKvvaU/F6P
PSZmsulFP4/ePH47xws74BXBR26+qtasN7winnmCq5+dDr289YGhYi+bvnsyTlO/
IbGSd9f1WAN8bi2l1o/4bX3lIwmhrdBSCeGIUXeE/HJuoHJgFgwD6LjCbtIHRHHM
IhMb5aE/QTo+rfilwFvo1U+DuBJOS8oZyf+jlbiUI1LI/D1aqZSNbGACkb9e9Lg7
rE5Nc77/29Sm7oiDn2w96DgLVXGPXMk+Z9ybZ/FhdBxEyWiqifvco6PMXBCIGjVL
2GTbLQKAbsH+MGKLKgXR7MtFlHtU06vad1QLI9hnKnDMfkaVdqGmJHRh2X8vNTyp
LJNEcWpzWA1Umh3axMtdVMtcgSIRdkVR/beXPwS9bX5Ecd+s8YUB3JTWcHHO1ed6
gFjMkIOaHtpxCj4PYcO9EcWKULb1mdGNp12i54tdsMyliN+PZLjYoxBCcFo+yIdF
ncKptrY0FdVc6t78Y+jyBU1774sjmEVlnbw3Ubciutv1gS040WWRg8zUPTtMNVW/
6n9mwHMSkT3PR2LzRMhegeTzs8+s8QCh9+EKegxm8lpn8vcfZqQrnQR75Mdp5mb1
OWsoc7NsvP3G6bRJNmOVgL9Z8Cw5GyyIxmRBhWscf7vfER6lIzTnPeeEzd5kexfp
Iw/6Yk1s8zUtkv+pq++gP4dp7qqrwY/mIK5w9vYZ6ZHfhpeFxpy5CjVv4HuTBSes
DimXbYwPkRXNdbmya9lcHggkYGEPJFTD13YULD5cO2C07e0cWPv8DinWFpvUO4al
zGTOGCWP8EV+cDq/sVdTC9lC+6SSnYhvN8OTP38nxZ+oy/orUzMvQlpbP6iJVBDQ
MvSRrATwP8csczW6Ywkvdjp2PR+KdQ0gMybjDq/IykjHvBlFTiWKxJID3EkY6F5f
8IqXpLtUoxiU4zXujp0RwRbW0FDjj8q+9jla0TejaiaSEvY5fwUccnsDsvLUBipU
gy+AUSEnfBWDkS0vhokiY8xZNvHQEj+fCZaiaF3vzmLVSQgYnozrlUhXs6rtX0bW
Pq0czINHQjOXoDwUqiFwKr+RLNIEjtpTEOLqOWz2skztOzU/0CWc8EAVjSYwPExO
3BTA6BQoGNyyQ1AGQ5U8jOB4XzFGLfygXsp1X7a+VcfhoNWCkHyPMmgxjoogCgv6
718rkxkoZI9e0/OfTlNEa8YtiYdiMA9saUReJLwXFu353QCD3pr+69KpIXl7z/4X
8gbRERKfDZJQbnE53EYlsBQrB477V7X3C7BJDJfbadMo55ULGCA1Uv8wax96Mou7
Ny+jQ63FF562fEjmSZVf3z0BtV/J7fOLkpCgpmDQ4xlNR7w1sDrIbjo6ELEKt95T
RQInHyyLKvsXftMsOFX8UGu5Wkh4iGo2P/rKPyZWkNv2PImvQIG51XZlEqdql2AS
WQ5v6jt6CBIkgy994By7QBXA+brITlxX4fQDGcob15Y1vLncrz9VSOGRRbLxq9Tu
BsAwPmBsxLcqOwDMnrW0qkQKQ7BBEvkB4y3OLVurxtxE95YoT+DU9gz3Nr4v3qBD
7R9E30NI8U+yAKHpGzdl0uloZgaEUr1yfwswqFKikb5mdneLDKdiCWjEhT4sIDqp
y0kHXpWwuV72CCt0H3Ttzda/v5VqCYJz5+1gIhhsxGpCrbJywfTZg7U+Jq7LNRXv
StnDlL1BqOXPbEHlffeegwARBlDS9JkPTlT9etycmvptxxMetJcxm3HrmDUXdFnA
SEwEpwQ3QKVqLVuviXV8Ph3FPZlBqq7pzDlKMkiecBAaHFUN7PopJKl40AycPwtr
hlSGFbyLs4oq9TSASZ7ZBn+MKcXGuG/cshv6Y0sVcnTxs7i4K8yWcVo8gWXjNUU5
thZxBORjHUQAnX9LFcTNh9F0VBSxrB7WqQXRHOjBU9T/HF/sNoVqJcb+sOe6Mkso
6GgJ8iJpJhKKvJ2MQJHokQE192VEuv5oohiVlfRYETH51j6bcknfIQggQUZNM/Vd
0Q13LenWrSGQzgcO3XJ2MViPa9cIGLWqct9LjXqo+WQB8CadOQh89jtuqBUtttvn
spCiGNoB0wZ+F+yFz4CztdX+O0VEOi8L/ePXWNMzWaIHHypcFhOa7LVVZ+QjEw29
4MK6dOvuQaiUjxwO6U784TSrOZt9yiwtQOvWhuZu5XzaifwsFxjxfp6ApY0hb3V3
/7CMVHzsy8LBa/ZUFG8rU42LfNXgJXLrdzqgSWYYSyQz64CkUecKyyKk0SsPP63a
jy6Dn3foRlTrnHHwbVl/t23mbsGyRUpGCT9d4W9PeQQbWl/3i2rHswqvPhKQi56y
8g7VKd9HMhpSM3M7NbXRqEJ9P3d+3OQpbzPZVOucuIw3nr8uM5VT2xpHeTHnyBqW
6gIv0d5cSbG1n6GIslJQA+fc8Z2DK7FWaIAeSRPlimCLL8mZvyVH3v4bXhXjHk02
9eHKKrIaLIMtZ9kFfXqf1uuQMeyi/du3ymQtlVjjA0bpGu3bdBlL169Eycg3DTg0
i9AcUPjMRGbN0w5lNo+Dk2+y3EUkjpwJ+Tjj5m1IILrGKzq5MHjo4f/9iF98XT1h
4bix7JAril3+2B8Rdeq91HuFzzfMdfP93gv9LghYa67rzgmTDxiEcWAzxgky/Rs2
DNnq0JNPIUsVuCZpZlT38TTs2eGA4C6/zdQ3QtkODJrjkJKt3c/tAU1Ph+i+8Dx1
5x8N5nE+UTIXefYyo7YObGrEe48nSZiF4syndbN8r5we2voLPblc8Eq2A4zm018x
wMIYB+J9bJw6JrlH9kYZzpkRALFLDlvHv5zDBRT05Ts0rIea2aSUnRBI+04I1d6h
Pvu7r38QHfA6h9MXUJayrrIAHPMO1GFVSiLujreAA6AcA+ZAzlCsRnH5xyRrRuV3
40rtq6vTNhdDxqeW30r5z5eh9DZGf1tPjU89loFyETY9BaljEVt9czTrRQE3loOB
d2jfm7jNBbglC4eFA/+Jf3W2Z2Tc4nWbRcnd20b17qXVPFZTPOEPkn/gJbrE+R61
9meRxXuRx941eLFONaA6si1aTC+g+8es2Cq1FXZzpyZcxjfPrsA69n/Ag+wuCNo3
mA4OPzgC7DrMKZP4+HpTCPbXWbtVlXXwP/RQkrJkM+zk7Mw+JQ5QuyGDsrfpzD4o
0yCQQVEMBeDAiAuRBmKFVWLpwIMH//n2fwKZGv5mSndmutjJJgPTUJCtiRW5oFYf
1xrRMKqzeonoQyzJZesY8ahgbttCeL/1axcSuRjPJxCHL5symhXrQWKpiAjmtl3E
TgtERtatFAjsF13NsicCMTVlsL2+Zv3kId4difq+6kJgS7q39mc81aU3VXJETwqf
DL2XTUnEFB2vLyD+Hx3LNZBE+Qss/VKIps3xG6P2oa9c4NwnDZWE23XTgS/N5Nu5
uYwC+f3SJR6PUQ+VQYixIW7PY2tIZoMRWM60lUCm5FeoFB9OjJNffS5+xmBJ0I6+
BtyFn2qguFac6AkQbdn53jvmZIfC8wh4wHSTaM1YxYss4Yd0jRKIWcZ8kfygwx36
CaGPsOcHz80ZdMZwADXbi/tw/RhcS/nygi2mBQV6XdbSKDYQzeD/C/Bxn5Yv4L73
Eg203oc3lEp+ypk3jbFnBkyuR3we0rI0nwD9TJt96f1ncSu3gRy4DatdWMdb6NBn
6WZrZuV7GdkG9/Q5yDkJXDwtHuLKck9YYuJFhrL3gw69tY8Oll6nRmSaG8zPBjuC
4pt9MgFV3O6tBPFbJyJcjoQrdVT6JyHOYF6yD3oD8i9Venr4ZcUBDCdyg4QaiH1i
u05p/p2uEOcvxGp50yHpGVHcLwN+rLb+uQdBpraNXSrVAn+HoWsKPDyfw1/lF/ly
mn9NkUZC9hiUd7S+cCYIhU4n7QvfQSz5onnvK0qK0OQ0k9h8BSCrBKU4m0UjXIzx
invKO67JkIC4cLlR2Dkv189kfFa6sdwPT+/3OlrxJxaDQ4YCh7pWlfMVeM1uouYr
TsUctSH2lfrfEAuEwcddN13WE/puEH3uxqPV1SPMLaWdkQh0hHhxXuaIB1LHAyTQ
WXlUSxgfqF5IA6q5EqrL+/ox/vzVEmJ7J9suoOHQsn+pGGF9yt/Dh+7kwpC0uxLB
Re05yiLh6K67thDyABE5TiEnP74aYyra6x8xvwTyxz0k4qftTdIw0/ONJrEiB04J
wM7hchekqPo0EuT0F3Rc5KNwd3HZofpphbdLvGkAcnAw+2EMLLUJ4F8O8qBFJCjF
VrLu95vU7BSOhzvesmwioVYjEKqgnPFNqkiarmITA4cNMsyh6j+35BD3qOROom23
gRwR9R+QgCSvhWhWniUGddDkXJq9G4PJDoGY19kbIJEqrNSCjas6FgfvxvtqCF53
gI8dfJIFs/dyFrjS/csDB0xVCPpJxmW8SiJvhI+hVB+AZJQ/iyD4RD6EYcNWge0s
en7JkRFJLbORfFPu8cMDJf56f3XUHTgNjIOi525aa9VLmm8b0821pir/03z8KMO3
RSCR9TF+Nt1WAiv9lR+Hecz0XGXnE+Wtq82ZlrKy8kEnKu/eOi1V1TteaYHJBEuo
g6FexOTRfk1JSI3xV2gxuTrtQRU2A7exa5ORzmBsCsk92miNKRX/GSaj/gOr/kP3
bTM4fIvb5Z4x/es2rCcKO90D5I5fXQpVt0r2u+gsR6VDfRCptKGHN0MobJE626eW
fOLEE205kzp6j1jqPu+xIigPvxTGQRBM8cD6G1pzZH+oq8eSrfI6KNPgxVi9Xe76
A51GxiRxwvkbSj8Qb2SbFw0O8jDHI1+PU+//N8AKL2hdVqzBQFz9vCurB0SFvaLJ
1sQzud8jDqAtrjHZvfCIkWWymh+PM5se/AcUe/X9ZZodX6YJomaOKIdpRC1Y26Rm
Yyf7qvVqznInJue0XrmIKcdKuVp6wUordLHiLQxzYsZ+vwbj4rIarBD+WPCC28BN
JVKxK2xB6Q9NR45nzcHVYShUwChHIQWa8+cRwJJSnbC3Gtsr6xJeD33jjUUz5vXO
LeK5BjqIRAZPWFTQuFsUNuMP0shnortswpL6pCj81Au283QEKItM79Ubc4Nr03uN
mcikBl97i9uWlWy31TGBHL7NxiYtdrTnY1X4S0T0B0w97VI7yll5wYVINqM4SiYp
0V8kZIPa3hJtgSzxOHDmoN81G6Nk+I8mzMwMSPEPpdcSQXKri/DUNZGaDzdyd3oI
+2jE5JKsZ8xisK+WjdoRtMfAYultnPtlL6B8l/sXDzDHSCZyXfLERb+CoDkurw6G
9QAOdvOw4baXxJ3M6RSCDAJi5M6afcQD2aN7Kwk2ldUfW8fTmfzgpXl03TrBip4W
QBKCSeMi80tYJXoLmhtGX22iE2d2BMXKe5A7nyHDDFPbkmrQghvjCn3q7/kDQqbx
sVjxelnWZejRG4lPCuZGf43ObP1mxl8SzpZtt/nh704Wz1l2juxt1ELSXPTR33Lf
Ham9ThAi2/KGQM74ANazjp7IGZLM8xGI3zjfBNHLCwO1Z0rD9BYsymFMeVCjAa0R
iYQtiQ+FzU8n/VRq33M8tAT4ULHQEunk0JBt8P6bUDY2RdB7RDN9SmYDJFKna8Xh
2H1UYUOzJpVSrfJRmTGY/GBOXDRgtM6JqiqsXsz0eCtxzG1VCZAo9/mEXZTYNEhi
Zv8vLG7mEulf/f5vn2HCZ02At7yrdFxl/tovAW4d3h/8KYLKNmOVdi6zKbjGtsv9
crfN4WsInfYlLdj+JMDtvSq+ajkvQD2xaxwsekzuSGjrIPTfYjAO51kfxY8ReS9f
s52uW5lDrXCRmMxD0F8lCrkhy+GUTv5SmB/87TAb7ZntHairTRIztxkaStLZXBhG
EbuZZIZtcfjCf2+8GpJw1Nf0sDXsbPRFWlhDfq3oMn/TEZJ/LLaQBBHCSSE4MmcM
Gc0Roze/DwZ9pyQHvZoir++FNU0Hr0v283LZm61OvZQaSKtnLSiw0b/IoLqGe0Rw
dqTEsrhybW/1ufqJbxdvUMeCEYIHbpRc5Cnf3EbSL7fD9DzMpL705qJrLIDzLCkb
jUzohoA/9NOaFhBH09H4SHCGT7H5X+28pbz/zT9Mnpy7i+vA8Ncp7Q3Bt29PBWDb
YTdIZKSk1KBi9DT0PMDAmvzfXZE+tr7Rs2WaaxNtsP7aGqoSuvQess6G19esIgV0
h5lH/pR5IrlaxZqCHc6E0J3dVEgTvlOtqsO12BtBEDd9Bv+GTBaeoxn2Jm4n5ikN
8PS587B7dB0Kz5ANeAMcD1ptXkM1Rqb/5qus94SdwMLMs6rrxoYBuqqeL7EooGss
qJYutOG/ezHSDX4G/EWvkj7K//TI6pSgZwo6U+Ti+DbvvPAadwqm/5GEPjTtlvcx
8rPqM7izlPmeD8a/IkN/QxKIlxvF8j2GUCnInEr38mL7Qb5++Hh0t23pQrUKxppH
iIdttFtlUlV1sLXXd+D1yH0aBMKgNyTPLPTj3ZjV16JotZZ+t8fRzty1Sy7OwKIx
ssi+chXOs/ZJja2bzYglLCsz8FEBgLr7V8MK735FDGVkp9gXb4fM1ayvPI38xN+b
KHvWvzxGzlzU5QsWiwkPo5+UVvs6WwEmEPt55F6hHftPAB4s8v7mi57bx+v3w8x5
WEz1b77euYpFu8SUYF/i6vAzRJclp18ia0TyH3HOgqzWC4SFAUUskN6vjvMkR677
Y0aIvxSwOKPInqo1rRWKd/qKC2+D5BPH+HRcZzf7DSlSjbhRlpCGNiI8gY0277bq
Ui8EbeChz3gcYfzyTsYrmjc49notxLGoDqP8zD2+BrHjvn6UN7M8l8q6AM0nKHHz
//3P258h3abb4zbh/jPVHZP4lpS46/kw0z7Bx07N3SQq7zbGnjVFLUfcU7nka08Y
odVYOdcvRZpXfhaSbxafHw1H0EnMzXHucnEEITXWrzsouPSOEo6lChDHzM66ksld
dncrboHxIyTPQ8Un2u9/oV58etgqiW+sEkeFEHowxUEyOi70QoL0wilbQ/zGG/uJ
2ZJS/VAcocS6QIzRHGMEF8Z15opgb/MiO15LOgQXPM4xWhqMvuMQpeYzm5vtrU3S
9JJH1gkQx1JAUdiXLgd8D5m63a9E+uxbisgamTbQUs0SfwgfKx+qOuGWxacQWu+A
colu03rAGNp0QqSkR/m54QY6EqUlMLdqqa+po8t9ypblDEkym6KeCF3mv8REI85g
R1lBHCn/ut8II5VqgE1fpPUwHS/E//5EccmeevyDIVpb3z7Sdqc1n5zGZKuVN2Am
yJnwz5uj6PnPOr3udFVxA2qV4TwiDVbr//nIF9mImpZeSYiYWSRVPeKkyYYwiqo/
dD22LXdqTyOrb5XIUCTk+3yrE1Z8Xh4mpqfmiQC75WPvaBi/kFQXlqz/XFK8WtbP
a4Kfq0cz7cWVybK6Q6t203rguXh+hzxKd8uMWiq7881qshq834A2EboNe0rHP322
RlVE5em6V9KAcezEgIBXzViCNLgwEtTjj/JyENPR8FUuuPjh021CWfe3q3zJu6ou
Msrr78xAA3fBaETfEDaL9Cgivp+FoAARs/tXqEHMgTYXgklvHsDRtpWPAPscJquf
kfx/ZHnqtNRvInEw4I4AsP2M/bumPEC2To386pDDOXMnMI0J0IKBdrdqjRbZoMQd
CPsMqxkiA3Ph31UjX9YNmJbh9GuOlNaRHHynkVnoDhw3HeNRiUJWji/sAKdoVibe
b0uVZe3+O86lHYIgafbYAZQ6+3K6wLOv8o+vbJ32qa1d0Dy69AoSvmtC934+PEZG
86iWAqQz6Pd5/JAuEFs2/8e9NDMAWel+ch1gCezHxA2KyS+meHZeoM1SFrLDczMf
RZRhjhNnW8nwPxRUdurL3jdyq0yjayItljuLZ9FgkUDCAYgJ9ikjTT5Q2vAb3AoX
oyV0Hxwkjd+0ezPOQ64K0dEErOkF22wUspb+wM68fcEX/ufHpWEa39p6t/OoIho3
XexIo3hTUONxxAKkOKImsPTf6KvJIeMLzMfVOK/op2lH8BJZyOiMQAn+ADOPJG9K
nVhfnjYbA18cUOCmgF+j3TCq+Si2KRgB+w2R+2/7m+bz9Q8Awlt8wt32JqPOqML4
KtJJKZgyYnE1ILXCkRS1ByOt3y0quWdxvcJMq/g2Wef+WBgDIOr615pbozpOk3OV
YJeUZoggj0sjYVk47RzFk2XFgvYzP9kfnk9GQahJF7RSyzLu4E2urM51DZpiO/uv
ncatwOqfOWrRDAMmiJLDO8c0LLC/LrgUF3nsGIUX4FeI79OIWsPWWIiSjKlFE6yv
w7fm7QpHU4qSGWGIWCEaz3OD7SEBoYoqwM0qMqfov7bBjW1KNwh0T/FVlZRjlNsF
9ns5fMk72jTX/OkDu9I6+80F74x288jP7Df1tMQI9ebE18I3m+A8VxGGkfTok0eh
bdzTWZXf9AiqNm7FTnuAW1vCb7FwzTo3bYb3LFn1DPkAjy1VdiaWOvXKByCf6vGS
mRBWUEyKaIR9zCSBVq3Es6djC0PsBTbFZFnjeHf98IpeqdLkDjma5v4hQ+XA9XTi
BcfaCEx+GQb8+GbUKUWWEFBZ63DKbv2W4DKJWUh+ehjXWoP3n3nLUbzAki3X1BDQ
ZeLgy/TELPcSbsOOJGjHQ5njoRu9hjyzFTO1E4WvpmrB3w8iOJoeZGuJn8NEblZj
cxW8XHl78yDwaSBl6w/4fYQKCxaL3HdFicHHhHjE47aqQIAyER9b5pOi/IcpYbPx
LXMMVrrmteOJ3sNbPt0TRZiYlEsNxlNYaa7l2mXyTCarYlmlxXXbkVHZWOh/79gN
k87ndA77eLYrk0nSlUYmhppsu7VbIWo53A5VQ1jB1uWj/UrD/SDrW1xkVxPanrH1
OLSoGKubW1DmIOmuU8dcc1BsrxK2HbO9WI1u0eMloqLEsqDUW/wxkiKO2OtsAHCe
+jgOk4L1KraPCi+pJdlt8kL7jumO6NBN0ysQc6hyhkqrudfG54++gHYeqdaLGl/O
41Hva1f5//Wh19pwV+JyfKp9bGFmPg5HPXPCmGI2MfP7k97bq1jODfJE1rKLMjSa
72c5RiuMFezkOSAZx8Ew60IlOPa8sCpbgQBmxiPngXOR2epChQOi3znWCLOFlift
ig56dffR1gPP56gVWLK+Btu8OmoKoHwdSTK4nE+U0wXtGuZmyqUKkLKTrmSG7ZOt
zEFx7rxOmA7G+AgtYGUuT4aUNcEmfczmlhAks3wRm1INc/7flf0icBInAHUtu3j+
1zxyv66XA9lW+BgCQzZpI4a9yduSBWU5vtpradlZ+4ED+IV1kZk3Fu04a56Q6dP1
/hNUT9DRnH26lVnoXQm1OBb91ef0V6Z80UZvtDO0tjBiBZ+yzRuv3TjdFgtGLTeK
bOJhHpnsb5Pe1fkvgYpUmSRQj0B4KGUP7KIRXn49XsYTCLM//ylAn7MDV5ti06Wv
tDWUMw+MYykfWK3Jb8otUZ4a06jJR8hkLYY8feV7ati0EN99Flqvb7fkBHFyQgn3
P15IoYrj3ZiGUunUEMz0ehb2tJbqMktQ2ypnNWsKXelqjg5UiBwhnnNAY40Qg3B7
QRec/twcPSXelAsUX5i+0Jfjkv2b6xD8BoIV3lk7w+t9LxysDGi5CLzf0jTYoyQk
nLuOtKhmvG24xJm9kZILFksR5I5VLo8Om3zqCpiv9erSKfpwlVzR2b6d7uPMsRij
Ti1NlezzB1KsJJrfKYAogBDcJfy7s4wrK3IS3KKCT2Vi2gHi6Ilf27RJBbSQ0VCo
VH2ct+pD+QErYj+53ZoS6vjqpivG7yxqPP5Zx3UsQnJFFMrbWqKQ0OGIKwkJsQCn
oD0lIwQf0+jXEg8efM+4H/otAqMvjNBWlxdNST2vVSOY3XaPt3t+Nlumxg/IpBfB
cTA8XB09YWS6IELr63heGHXTHJs5MwGDZ1NbpUZcnq2DxgSA9ViyF27M/0M4XJkT
XOj6WHwW13wOPLSrMVmf2hViGYLw2nkai3IXF2k6fi+Rv4mCN76h8L4jQ4pkRugY
diOD0DKtLYkdH9LIUAEfe2mPV6Vw3/hHL6FOoDXVIbxadqWA1ZIJkXqp5sX1OoXD
owVxMD65NVF106sWgSKIbxrrsuM9Xy0P4BjiMaVAerbYSV3h+Ss67DwrzLKruc0I
yTHivinX2Yy9UslXCKCTx9OuwV1nOHZUim4SMSxkF4ug0izYjR2K/SP7LYOk2m8P
cGcJ/Pei94uIU7yEl1Dn+Hfadtxdd0dh3E9RO1oDSr1NHp5VP0AlygjS1FIP54A4
r+9FuGg0KKzRV9nWDvfkCcK/Kn2TOLK+9BU6o0AbkybW+6VYjK03CmH50iIdlg5D
A9SSQwGwtWwdr3hRAu04SD0qzQJ83E9WWrFQJ0qxBgKT0HmYsYPuDyDUhM6BvErM
xa66djuHhIJuTRzKDZssbaHMNhEjFd3gNe5cGimj6hNiamSM4DXeGc8VOL6/2YDt
mJP2YZp5MPvFRxCBO4S2S0mgUqodG/nT0MLyn3BikDYSTE68Rnun4AWY7RBlVbIX
qOf04Sg9TP7g+io4do8kfnQj6E/CvSl5P+CgYxYYV2ZmGqn/35uZDc7yVtpfF8th
zPLuUI1RL3RF/VheqEgqme97vRCCJPFW9UkR4Uyho3y+utN2bhZKRvOm84ZcJAa7
nUnKfRD00LCRXCGOdRESrC5DlsneolyUX7Zt7MdnU1P66VJsf8HtlGcrjqEcox5N
KukxinuNh7Oixkt6Zo4Ea7/xkGtU4Ag7w6NoQIgKbGwI16X66U8QL0MBq1XMOltm
/ICrGIrCk99IenVpUOcDd6T+/msKmpDzZi1w4LLu43V/FEdCEoYYb2oXnYnaRuVb
bzk3pzHEReRu13JLKf/XJ3fdN/P+bPEdhbup1fWqRzfGwSIr7ovpf3QL2Ukol0Rt
VynF5fKr/b1Csv8clj/ToMpPCrmwjAcB+AzhJ5jfvtsskYSYSWi19lE4LbOjSiXf
bcBl0BphDCE8pSVgjlphoNxJm4n6tn8rOapFcrYfylnGsGqmVatrg4ZLRGvyAbai
3QzX7eH7JqauULOjWE/84LXwpjFiLBf6+u4HDB5gZmJwD+6LnkoQtDFVhB1pBNw6
IjxPujKKWytHNMi6jII1VoU66rIUZcILKlEpDhIZlUr1zGlsKDhLkwGNvBkIuIrl
S+nrwtQ22pGQJDwRsSAUQqtOumFt/Kycn2oX2tdsbloLKOSgarSY2xWdu/xqh4E+
oZp4V10WWG4Tyu4oPNhu6ek6uySgDR59fBYuPOHqh09N+x/rgQ9Qao9/IQwIBpu9
6yahF4Ty+Cp6djY0pBcqtgsPvGrwj/psvhtat8v3wMXZg9Bq54tMAT3occym2bCo
sNCJSHTf9ds4Yz+cG0hHe6BB1nhiSHCgWU84RIiHDM6EdI4TEgvTgU9QFNA0Zo2u
h/baVpM1FHzFJXIZ4uJEoSA/RSy22oKc2cdwkFCraY2bMfWmQdql1Hi/QCiCmjgq
xEQ0BoxYjBivX9YC/L3m/7K4nUnKh/12i6lolLVCyFd0RtezU/wLX9tPGZq3GUbB
qFHeAY4euKkrvscAEylSWbsI9ceaAdQd9u5DnbuTEmeqL5spiFUUmb8Qf8VMqat3
a+5W3Y9TBflu+Zxz7/1gfNkd+/FEWj8YtWAd7ENWYVN9H5VOBOFrwIGSrCLEMG5B
lWcuE3sT9XGiaHAMk7F2nHKfHnu3d481icJxPejYeZLuJaFxv4qwtHd9DNggLUfa
z/SeE1WL0mww31iIOu2yDRNbfTmeHbB6523QIirv0zX7i8Q8IvM1gzBbT7CPA7Vf
3MkrBtZPsQgEuLzkDjhquv1j2tMn77dopzucNgEu50EnMaml2dcOQDwZIfnAFT/Y
K70GTiKs/7MRdwdkQeJRl9Xo6ul9y24UlX1DddNxSWV8vPqeNZWRQXQBo9s51qkT
DyLVhCCJ0vLas7O5hLMJc69XPgFdHThov7VYgHY59y4oTcvv2vbvfGR7kCi2XFN4
3h4tVCTvdDp55oimucscd/V1n+yclIjuSoc3r0lgX/16if1ObfxiOTRCQrMyivgN
61bCaubOwF+SR9BWB7r8TS91wAMi6jw0wgw/4kw78J5Ee1VHBsFB/P1eu+AH3CbX
U9bGK4PEmg91byorVdnW5u1EqXXmfK3RjRbwCbSsgHExKoxrr2bSY9IV8JcjNts/
8w8/ToZVVhaykDin5Dut3tyg1h0CarQuRUkX9jBM39C/Fm+Nll8CCt8JHZ01NM+U
Kh3HFHOPl/xwusV/qg4UmnJMgO1yoWMyK9vqHPJQFTZxOtgFg1Da9lB1hSB9oIyW
T2jBJuEVuZz4/abvOJPkbLM5yKClviUkxhphIE4ORWPseq5wnDTkkaZGqPIX5hgb
mT/eVkciDUWfn5pFaeSoe4YYS+l50KEwlikdMxg8vevJeJnSp1Szq92wUH/yMCuN
QO/gT6Ylm/vdOpbgo40xXHyC9soR6bYV5Lk6ydhZTbRI7A/6P+ZJ86mKB+YxCff9
JsS6QpAS+wAETD7Pensmc8YB7SSEGyjX52m0Mh9IDgrlzegLevQcaLiirYQDV+dP
ApPt/tH9nXMrxmvX3YtntTYnLGWJErswW3mL0Fu0YtarPLhSqfzKW5piKRvRDjN0
kIW5JhPD6ayqH+rgzubkAM1jWr1BQ710N5EO8PcBwpJ22d5jd3wzRIvFLX5Q14NO
o+mrPgRlU/8EPOFvwktMCaVuFJsnj3mg8lkCJgfVaZ8lQuXT2ToB6WOWrE4Ywspo
gvfEC7hXxZHLInUw4YlIA3WXawc4qG9bijdog4PJhdtmtI2Q5f9HioRzp2FBJd36
MEjX3W1mTHDoz2uU1TZOVOy7W/ML7K5cviZa73Q8Ru2gtSQhomO+rcDhvFCp08wC
V2V9AHFRjx4qA0cfQwEzO5cI3WFbh4MMr7eg07rJNxESjDqt57njMZtB3Fg8KSRU
PWuzPpxvqbgqWXuv8Dk03Z2wJyRJj6Sj3m301AkR2voU/vyt+4j0M/GVX105kqcq
pm6EYfZOxDU+e/oSrgqnaEmqV/BkwA7ZlCCGgqS/U/YfZTdiX+ImmP4UE+m3oXOs
76GVQbO0qJlAWLnvWLP5InLOJxvJddGdy9TvZmugQu77qnyD6RO2VSMvVLNCnjLo
uEaB4JffYAxPIVPq5ObpejjpMFFREKPgmfw3tEla5RN8vFiwYft4+4HTVIVnhuZm
/Y7eLRKO2ai0LeyD5crjAfJOyMzHWhC/k8zGzNn4OkKVDf4czw5rFYYO1WjZKJ1o
NQ92RX9mybma7c+ooDUr9NFNz4rwVOnyoD9ZX9C6IKjgxk6Q+SUrvtDWEtKLpyDk
9jQRFNKpZjP1UhUyXSy4MmttWAe9Wa0KjOIvmBRjcD8G0/Leq7f2ulbvZALNm5Jm
ELplHxt+Toe/PhY+0T6b54ykFp4ZrVl4jEKNAfkslQxL4umhNPEc9fWSAbx9xHhf
Y5BdQNt9iRxWdMjR4NWeMzZVzSDcL89oJczo1Awz6BhFDk6RiUNuRN++Ms7pA/uU
JAGNQ/twSWjYtIoTIj1eYIGpd2oMWl1pagVvCua7+emm6YG7UiVvd5Z11HgUlvfo
5wdt+o/dJnCwYAKLVMfWs2R5BW2+Ng8uTlfqkCDVcuc+p08nnFylRUmJa27JrBKE
Kz3NDkZ9jK1w+Nq9CodPriWoqn6+KjQGg/VnWv6y7OZCbYBrN7E1ZMXmr57hZXYj
JwRpR7+cjVY2yX7LQg5Psxdw4pBRfTB3HoZpcYWZAVRg0X9RQqcZ/7caEdCs/eZg
PC0n5GrzJzzIsLrPbogEsq0xtkyy+TrQ/Hf0n1JKbzsuGv0feQ73cOvDOXpG1+s+
AXcvKt7YzRZh85hvJvK55DTB+W/QK63LKcb09Tgu/gBB1H8dWpgqvdZkmNawkiPc
Z3weQHDkMIcth0VOjwRk5y0AwZfXjycF83R4tls36z3kP2L+aTcKb1IJ30jWDo3g
LEqGjibouIA72n1oqO3K3812zJoRbz0EKtedvwMFAms+NqmIE06nI39UaiHORPRv
JE3eUv9HkR67V3/gJD37724j2gIXIMzxIK5vSczwtUcJ8IU0J3DFfmysaxsU951i
YFzvK9x+ncxj293U3Ejt2myvYSsbWQzWyvOLEmjlXMI5bWucycfFwDSgDzfC6j2v
IBOqr+N+K8vptyBWQelbmyV0iENZl/DqmL0p74zlP5afHz/Rm2SCVI0E3jQdciP5
NNAk0/tn3gXKL4T49Gwv6DCDUoatPXxb48IquSn4rrabXS8gmymJqDy0fFthhfX+
Prr55BpKvosFdliIIcvlXnIHIW7P2siTyOPf6E/bYty416OlZCcFhF/Bkql/RT7h
MidQ7KeL2JSsMfChSqhlaDOtxGvsr5GDyQlM7DUkJpzgtqghzwvltj9FzZj1P2Vz
112TS+SV1O2Gy1rRa4ke1uWIDOHAtXYqk1gbrTZjACErbrkBhDlktqk4gh3FWVde
78xf4/2jSw2h87E41aByCxuVOiOZW9XooiKJpVSzT2oGSrR94TfY+DdKMCqQntxD
uelk21tlQaomFk7N6KKipkEG8e+dYNbjyafEUlEsrS3XlhUPgGbPDT/Xz3RIovyS
hygdIbJ+prAo+abKRU/0lzTUIerSbmm0YUWCQPqca9HW9YF06Ytwt8ZCnJAME1ae
EwZIZlN+fT5bbziNiDRxFSuWzMeYwIe9ijJtlm4K804KpEI+RJhPW9jAdYmnk8n9
+SQQmbUPJMqIST9ICXQ4ll3KFg+TGsvQglCWmTPSrUawLMNbGf4ZW362owsF4IYt
W92qOaqQOEIfaZXJLtE+q4v66f4MYZbfd5tJ6+WOXi+Uh3vCICe2ezZUQLfreTC6
gf+5QggHLb2rIwNTBghp+BudqTvlw+/JYIgzNXt/ogambg6IGue1QsjMBfPHYAA/
WGqLe33Pl0JO+BrheR0ih51JXXQ9kf9VN+qI5WzxwS7DGOFByF5f/3anVTdtzyRn
x/YPlAPWjx0nLXCgtSmiiE+TDHBwNAtg8M9cIHvI8v+PVQw7h8yAAP5mPEvYZ1rF
mQmUEOr+i5Ev9G/e0OwpZk8SOag4TPqMQbYTt7YIfCd2EHg2GvwbhlwTv2iZfXYk
x/eRqvL6GWsYHnMPj79agpSjvijlEqDVecJKuObh3L4GxQibE0no50VF+EsolQQH
CAG+z0sWR4Ya6lwopYKm+LQ/2jdRQxlWHYvCNUzq+d48vrs4xuOYr7pZ2dZfM25T
XNsGoboE3/zuxP5Pa4VeWeg1glf1haAvX0l+oJg2YgKL82ZQF6X4T+8OA3/OGi4J
8SBHq15pr+8zD3l7wRe144kUdvQ6ZrTsssN50AfUwbyd3w0Gs3NXh/77V+f26/Bx
yixFnq1lD5NxETK9LqxY4gsJacA/cobvxY3snPKwL9BGcCna4NtqmbK0qQKQ8DIB
GiojzXuzJPaB1P6mFqNt/VP7D1BN17VpvxzwV8fvSXyb3DKN0FD2H0txa0m+Wz/M
ynK7JcHtYGjFgK9bQ6uGh4ccZ8Ctn3VM3AWUBR3Vnww3NliYL3NEoJIJZdnWvE1U
qbrWyXHbuSJ2QvbqzYsUxjPZ09f5In3rqdWHMrMq/pjWpWBk+SO793VudNqa+eeb
lQVUONjYjqPc1ZcyjcUzW+9NNelA6q+nZ7nRWJvfz8ADJu4QVuCzDoykE6TdFOMF
Lmf+vlmlEQ5ox9934v/QBVghrGIxLqjHSiPKL5s0wBB/A6SD1jgm3lK63nf8lK57
TLwyn3CZwtSovmH9yikqzxahpECYEklxbPn2QBfVTGynz7UA+cY1EG8gnaWqlF6P
+DB5FUysvi37Z1aSgunZeJcYUDcu69C9xPXGN6AIap5QO3M+OuUxxaN1JYhZg0N2
ld268JdfvTumtUjDu+ZeKhgbgdzO0RffRiG+gBAktlmluptgvSiaMlpc2VJunxB3
yCOP/OBD3T27z3mN08SwmfRJAqZd4Dpf0yyPhUftfa86TwQF/bjyCoL5vQZZAAG2
7/SYCk4pxbHjRSWnvX3RdoKIHEaggtQcYRi5hV2Id9cPSwhszqDRPkXCaYyIOChi
1qPCT4zyb7OsUaBs+yLbDgv4t1oMhZ/PS8vdL5QfTjfX7OOHZ3+1iWzr4yfFnxFI
wmMYnfVwStuQ2PUuGEI5Ys8V3tYHUPz2LLMeQcbqIGmZuOYXugMDG8L2om+GY1sQ
6rxHFZ9Ft8GKcHzszRcu7Fvlfw+SLwmjDkwoSyU9dYKaodEAKRTfAnEAUXyocBvN
e2i0ddsam975LWV6qyduo+PCIgeLB6ZShHCiojeeiM/rDjDtuFxLnIWMpEJ28xyN
OJbWrELScfnmA4LzlDNrOca/Rf1yIK4O0jghDlla04vnZ18x+txXmYxIr2jotfqS
EmLbopH/E3I5mi0T85hHJlYWsrGnS8FWgY4RpXhy8e9MPkiXhurwIl6TOrRRGr94
yxvJ3RHEEIPbltld+EY3jMU+VksWRvclSLb4o8hMDRLLxMLQQ5fFPun7uLwRtsvT
v+zQE0bADS8mHZ1w2bBzhq244gKJHxKuEfmRZSQ7r7+B7OgDbb2befsWy+A0W9ny
84xwShUuHmH3NEenJqr0ohZGKf18w/q9vhZipB03aATAu2nD0mQyPAHgvknl0efQ
ph86mSLB2bqBy/SNen70bdAlS8bc/pe335ZQ81j/yaqCVyXjRrbXd9XizWW3Szt2
g4hqmkDWJkm/R8zVCm5zZOHDpA5rl1rAWz8nj9OQHCe8bBs7UR/7qd1djdIR2ooB
PFrgwOjMZ9anjezh1Qy8SChbYeU1tVu5fP/EyjNsRlBJzOixDqtOikfvOYrV8K72
lMLt4709VVzzmHIce33zMxmW3LS463dZxpA990Lgo6QYfOcXxm48ztYWId153ZZX
bDTGAOCcjAnVOF71ulNd01LcBzOJX8t/e6gENnX1fpgMky+afkWhovSryChRVotJ
j4z0YsjGPzliFG8m2HgftJ0mPr0vqa53TaPSAzlo/5+AjSIGoo169pJNuHnlhvAD
koAHWY3cnoM67/ezehbqfJLyonSauGbLyHog/QI/JUBxAUSbQgDeamGEYlU7prrF
t7nOE/GVu0Xk/P0S1fJIhCF7hnk3rcgO16gb44c9PLh98jUdxV3QoFT+jN0ldULF
13a6lvNvz0WQzMozt3kHcIIqGH1uYEAKzC6ahru+mDEpxSBDtis5dir/+GL7A+Bi
Dk76n7ULHFYZJ6fa3MTVA8Ej4/3jlpvQnukxBNz9pYpU/09EgzV31xnlIX/A9c/w
Vygwm2zmETRVsi9BQBwkK2/OcJAXY8giKHcPFbC4Rzgq6/H45I2sG0Kj5ZrHdgzv
uB1+VqzUsGntK0OE1mmoeneV04FYQuooV3idcy6QYh5QHa5Y44+2nTAqs55V3QEl
wWFubO79QSRSzVJC8dfZ4QgeGvsiuKL2T2fhsdvFT8cyt5pIc8spRsWKfc/yLlo3
7mR7fuYEc7X7n1Pk0MvBQ7NL9yRQFZcosMAoHfDj+ehKlCJumU4lGu8D8E72YRhw
hQpQf0BeX7UimWvHetHjTqCwobWyVBKSIhDZZtF+EOCM8uQpdgIDLvUed8CJE/NO
GDEcyKGzu7Sjp2M60RniprrLTO+LQdbkEhTj76sO5GlmutCLuWw2+Mg1sh3XTAiY
Ui6I5KxaeVjtp6BUBZCUophjJXK42Blwydlx5mwyvL2IMQ4KMo447pyA0LwAkZQM
Eo4zWzwO7LxzYeo8zim+7bmL6eNjXQoftCg7HB3xjfstgjnoX8DyAX80yKF4AI45
gFLd7lKXGZMXNQ3AwlQ/gpe0OIyhRrQnH4htfezlX1D0HVSnThss9k87j/Maa1LQ
6jczFkCm1Omn5uKogLj1SWKn7XxTkZPpQQN1XsdB/+zioe3ld0/12A+ufQdtudVx
riBLb23WFIg/wUwGfHoPsCim3NoRMuOqiuLS+efRXeLWZNCcLd47lG4aj7OzjL22
K05YmUsp7s8dfz5qu17uzs+NDTrsRGKpQym9tsxPeEDE+YTezxvs8MqGZrKbojQY
zV//lVg6upAX2H+4LaWNLRfMaR9tbqO185TU4hFELvjtgYBU13d9Umb6/GLwACxI
4WSk7kK1uR6WQCD9S5/YtoT0PuwGZ2k1l6i+9A4PvT33bdrJA5D/GEQByauZvoWp
Kewj/K4ZuY7C1fsIesBACVuQNsuf7Wl1gLBmP4RH7tRXoYFAtWX0LR6LifkpFtjW
19FLlmCwyC7fCqdbv1RmzsSpWzRaTD+U4JmUShYLaTHsurFi9RbGcoMvCvaHJsDf
6WZk0Y1wHEy/qOSl/VxKiaHPwdDN6ZvnEaUwxQVRn2M+7tzE16JNtsAdccQoxc5B
aqTc4Qhz/ZBO/ZtWLuKAlR6+WAcvRKzW1eFsdBFInd29N5ZWfyXhNwdG/Pu/O23d
egJcFJXoQLiRF4cwN/SZv7CJWO5M3tB0i0NkQs1klKC86fiwAkF7Rg7o7IEfXt1v
9zUMl5RcLBJSnAEUMZR2u88SMTPtOGtrOjIo+NOm9hZhubWDECKIItqLTAMJGS9A
j3x2CpUWX9vorYH1/HCh1CSLXL8tSqIkrGl0b6x8kEFXumhqKnlDULbpCZ72UFJ/
qZgEyCZuudR/sb+asc7etN88z+NUggiPu19jBLyBjWM0IezKDgsgSa/GQ+USV8u1
8q+0fyrEo1JDby7+KqKGVK3RM5KudbpBOCK/RK7DpfzIu/Ikaptiiq8KK3i7Bf2U
bN/Y5NNzWGtY80yUJlJcTGssYe95ETcRFXXI7fyCHpwWnshtuaPSLN1kPKSGrpSL
Yks90XWmIjfy2HAmUjiljCNj142/ZtCaS69tAe7SdYGA6H3W9oLdPNPWyT6r3hdG
ntFT9yQ9P972tFb6w2TIswutxa6URlFZ2i+VoncYy3l2od700vIziyjPsILMjrT5
aMCG3iWL2WYA1KNEBlQLY8qTQGSGYRDt5Eu3/AbHHo4Lw7b4GvrLt6QLL0R9o29j
JwXhmZ3YAOVbtqbtVr9Duumk35W/p+R3TAEiWnj5bugww5qqRCMEJTt81tqSLtzO
C0ov9z8jgJu6W4d+N+z8JAOGadTQ8Y/euItv26C4OSPJmeGtRFpcrmarQDXh2lfV
enO0ey5r6kHWCFG67iWe+0nVPI2hwb1iE7UnRjYPkSswoq6NUSzdSUiOlKk0aIXm
cj6RNWSGtxAyUoBUzAEOvG3mYnC9JU7ykT3243a8cqE4PRCZAx9AO17BXuuVeLVk
iQUx9Xx7BgHMrymd8n7SBddOPAPq0rmkkfD2+qLtPBV4x49m09t9/ZcDSWxLfAXG
7TinFQRe4XhMlpBKZIteB3LAnbgHsrrdyD+ABV7QW28SSy4NIpcZy1XTVF13V1Ys
kgydui77pB9oZOBNxu5JnGQTD0tArLwCj/mrRc+ohAV90iIH66tCoXEqKER3M8aG
v5VE6N7fsDsln7PdnvPOVOygKNN43WRA4V/3aLrHbtxJk0IpNBZfY4LyL/yghpWx
KB3b1rfkzN3rRZG9i1+kPUGp3tqDnC1DBjamSANySzdykfQgKlaYjAD0NbfLolsW
MNnRQ1uf31QoAYdRQT3fvSsg6ND17hi8B3X/6ejoYduZiI4QM5RsIUoMtcoVvHQK
L9kpBmEvm4yQnBxSCl9YLFJWyV9En83wQYPVBrj6Wj3Y//ZKDsyWP5cg83B8jna1
gWmH24GD82HnANbCaNKXRLqnEucn2rsIFhukhWhXyLGrNcxaOqrCneCrepYfe9G+
FulploTGl1oLZGfeiNmEe0x3SjKKBKm3s5iw/xJx2bl5/LWRdHeS3VRm7Ibi3rAk
8EoZe/qrWW2LVkknrcscB2EBpQwb0feb7H53QiR/8Lhus9jCYxYPhK/LLTpvKjhP
3hBvMMxTUBCkKk9TPx415BzsnaPqaOk6LVjs6Cyysxs5voDOZfmTvCPn5xKs+r8x
Zg9zpCIJ8YkC6wBn3YdQVtTl1J/XH+QOtNOXJOTN0dtJ7K9R2Ua0YyfnzNED/9CT
t3+UnvOFFxueE7TVB/TMgRrYuzuK/LCVzhti2lQMFDlo89UZXNMq/2RdLLwdCSoW
0yd6drDr44KKy5efmtAv0xjqqQ7QZwwaFk1aHQM2+kmC8nQuZQW5ZvycT8QFFbFr
lyDegphIOvjsQx7C3t9M43CC5BbnebDKAusU1RZz2TVyzWmFH0YApdvvBxTHCshw
zL2IE7wo75jXq3hyQ6+X5V795gnUx1mam4/WGf3Geon6iiOL/jWmrIzS7JshTc/k
UCaT6i5YxmKQRJYR8xY0ARJ6CLEriQlSO6MaYlFoUJNQdsAAVaIWWjyoph8dAV+S
m/EyZqJCisjKQd2Tyovvk+O1oC6lzzCp4RFhVgnhqID2UjtoNcUzLoEgG4S7LW/J
tjkiGmklBNWi68Zw8ZywWpU0cDIyM2jtlbpJZyfNCuANP1wca/E/YzUSkNOF3m90
BdNaBzZGt65uNWzVAna/iuQyW5f6AWLlLafhHgZEDFDC+dSFwcyvsV7nRnYsh2xF
frpku6CCmc+7pSlV8ZUqMnhf2UqHgSGApsl+fIPHmHaLEvnJqlgyIfkz29p4avnn
NosIgtIZ88IzXYDhQkf44j/SQrZ7AIYB4pTrh1W/fIc1Eyj3m4mY/zogmAsBImpt
8JjbtCBFZUbqiUzH20wKA5SJ0nRjnNObz3B/9741pgwen6YcuUKqjCyDhN8clGtB
J8PQDSwGDdWMijeV1s1nsA0w5//rFlT37TFOFC+NKeMIpFa8Xnfgpf3aRQAyB4P8
lr6akBRs7kq7nBDGs1Q/0c5NrmIGcejk9pv47xqJ7vMt7mRCLuP6FnnOVy9WXnFE
xBsP1QmONsdx1OJi+cpXCgyF33w7pZXRBOSU+ksgmlHBgDuAdhS9jJ2GlmM8XzLP
+g1beo2jn2+yqH/OhBuVTW5rPocvvspDi4f8LXoVaCPqi/ekT61XP5VLYDu3+7zc
/8tysYf0zoC/RaOw4HLNnCH078FZCSD3uSIuVM9w73ovsEJt8rWaU95f4zV1INf8
/Yy3kNs2kcfHhVSs8kl5fvKuEY0UGgzappbpM2N0e+6num+eN+hxJ7ZMNAn6i/qD
2GI1ccXGp8Yt5zHg5J+MgVgZDIKOBvFj62iyYcQfHg6+Qi6dZeAFz/RU7Q59jGss
rtuoZxaEsxj3RXLCyqYuuzWCdrqmi8hkERKaWVuIMhLdphqyJ1KwMEXbmQ8ErWII
kMsQHRyP4xs9oGv3JMnpkGcHccd/wkAaJ/e4njmBhhBAc+iOp7lWTL5tWFYKWm+u
eCw2X3kz+rZYJSih6ozeVAli8B81+ySb+/tqON/qOYM5KrwDKsxOElYurzm/YRZG
yxq61OY+Kc/KAdEbVCBI//njccueFjLOSgyXU97LYpdpHb3M3h0bjsBScO1qBwoQ
szGrTYmtqzfDdwzXHCdJNSJn8rTep8Dbu5GQcy1+8QuIPwT8ifSmpInOo8w89tLx
hnkROTQlC8bUnZVqXBRgxphosYH1+LkdTyCmvHMvb+1c2IqUP1DkbShy2gPjBfOi
d0iZTLFwjR4+Oq5p+sX96i/FxdIoSbYJF5GiNjNhGKj5q5fqMCCISKTs3ICKcIrX
hdDj4RE/gYLQNgH8cjOLiHxk38vQT+XLHn6tGOwnNrD42/+BjT/IvEqjc4AnnBvd
/2wC6psmbkrmXYe/1/sBukPHUnaDH7oviLtcbTGdSSuWqzG40LdS04COMooJV1Kc
UPK5G3UPucK5moQqlNKyrYqccN5Lb8zHvFqZ6I3dwsx+iGDK+Ky9vsLT/DVsTLgN
cBvZDNVpyH3AoGViywHd+iw4M+rwOy0NRQbCtxYejozLXhVeD1A1pVHR40Pae461
BQiLCjBbdT4zzss05mek7CUveJBjpS6Cq3aOzF9fLSa019mQCMOnpG09C+ZkRiNx
jAyBsNLP6ioS7pQAGGT1UyDG3ZI9Rj+7RxIFqy1WAeB3ywktlxoXLzvEyZnekY40
CcflMWHweB2U3jUw36mcg+QJDk+S9Ukp1fauAaJc+jQLoSrjglxqDEbKdEI1uafm
NK6vDHuQjQxQhGrp5QRPX4oA+BpaxmfKX1o4Cn+Iw4eOe5Jv5dOM8ueEi5CwaEi2
VfobCd2lCA0oO5NCSChmVJGjlWjgSzln+wWDYLibO1UIR1TMPcv3rCFgI9sqBsLi
XUM0m4XnEsx/bxPRP8Uf2ct8N3AwlUsTWkbSSp1/K/DOYcs0f+VWl4qcAY9lMVsX
HDE655ytQe3SHlFWuDVBwyDhTfuF+dsBZ+gITivCL7HHmJpJxlAfSoyhg2tG2W69
8AKvIHxKN4De/YRbbvL/y/miaE5/0KN00bsFCJWw/1SN00Kk7a1vxd38LnfTuWwT
bj+KTxjOtkj5ebKscP945LdaXbdxWNWjG3uo0ELb8obCagRGsb/ZyXRkWibkNfnm
U9vtwjYTH9+ib7Q1lPzDgunVsjlwfha7yimTJ30+qrZK7LYALmI+nlKKVa1sE+SM
VsbVpzEhJC7HP0m1K00lovT2awfgYAjLcH9Ozhk9tU+J9gAIbvZ47MSSBILT7y4L
iaMUSJFGC91I5B3P5LxWIhOOGf+PGq7J2ZNYFqIhDCIXAuYmW6kGH8s8mVii9RYX
h5Nb1HcfrknA8Kz9qHNI9DjxtuU1AJ77bDVU2l+GQKtxaW4wTeW2qOI61Ysob/hI
Bb+I9+wBIGYi0Mx2DiJvEFSxfYwiBKgy7qwx7C5zbKlLYBzu/yHaypHOisa1JVFn
VxsdibIBE9fEvUBFypDj0x7uHsGvqjU2KblF2a3+1rwEEx3cbLTCPU6ht5mnTHCJ
9bgVDAbFbk18657yGqCpwRTlC46wfuCm/R/7GubjVuNq545jkWyH0hro2wiqmdnb
OBXHTfVhu0OLP5fdhUdPkpMlm8fHlQapn+7XTAlBqECrdzlRFxqmQdnZB8fCKUMH
ZrNbs3L9Fc1Ii/P1hlS3TufQ/s6drc+HeSE2ctx3T/SoxcZ8AJCq8ooyF6Utkga0
A8axFx4XdTvz/in7wWzkgxtk5kxhWBke5yIPtO4vwBm0jytdPjObaKvQNc0GM3Ha
S1pPRZu6dHJVl+osXC01W/7nSZZjMjTiRUuaCNF91AsW7L+Efn4johgMyua13cfC
QX+jZrEmm+ol07X1CAh0MQTog+vITcKilw7dLS+MWl1bSdx0iGH+L516MVq5LEp8
7/fMQ25ecY0BzzPWYIrxHl52y7oYLEoSMgh8HBBT1P269VUo8W+CAxYsUCzN1Qz+
hRqifyXoJyIcMjnHee9rHrYH3aG1PHb9FQObNDxMHJPBdfbAKUXsR4DgWsTBgFEQ
YBiuV3MNvnfQ+FXNPGIbx6sNMHXOHLfngDh+CDZtqHH+bGTEngaoV7npwQ9jAymc
j1OiIgY5UUw4Oz24cwDpKx7AQDrsV0hUxBWYLBqXTKOCffvEtgDSyOztiN80WAeX
evEcfr4pTAP2E75Ku/+/ng8gA/9qhJo0xk+c4c6ESOBLIPgJSLwy3gePxeTaEwKk
sGAT7r7TQzVW1nH6vu2kX1j3ZNUe0WwUi+Pvw9pbKva8GFSc+W2T7d/6PEucy9UG
AnoVgNYubY/JtYcvZFvvR0xwraTTTy9v331Xp1cyWeES2oAaMmbH49S8DW5LE3o/
LGLT2yvxQQBjhhb3q16twOote/C/0zep6mkg4rGMKW4X/dkVTTnqy41ziZxudZNY
felXBrzUwUiSToOHFP+JlMPDKRvp4yzAurHvYtPT2rYoxXzmgKEOY5OEDwWUXuK7
ASZvnXCKLLsQnbNN7YBxJ8fu18p7U2NYlUi99II1n7oo/fO8o2HHqTOXBCYpHd7Z
fMRFA8JwOntj8oy2Y0uwi1K9jkqxov58+qDWhs/dNWeRkibst0+/UPNuJ/r6oUUa
+2oygDlLNR7K6iHdW+XTobQEppOC/QIc6jlovIALXksL7j0yPzV+H5edeSqBvABw
c0rDMtO4soVLeAXK4xwuLFTNiKCIoq18oPnxeBKcCG38+TxiE1HqHGuQq5yb+nxx
+W2QGfcU7eWELKt5jo+Auu5jHZyWf8ga8BSHL6/6QVRzsHw0gnDbmHl36J4wZ02D
Hd6F/HQafr5n5UGJZmvxqtpGLJoVcT8Kp2tCl8PSu8dF0i1O/IUyG/b17ahpZwYh
i+xkQ90OKf0TanfQ8DCNg9mzwiqZd5rU6Po4fXcvBz2Qel92mgJc/mK5dayIris1
tMMDks9XpO/2isVMQYRk7oCujvofL2aKngCw7VoEwsl81hCPg43tpN5YHgHqwbWa
Y0s0BNzdgiPQbE7VL/eWIx/N4+zQ7jTewUcna0XMOYDJjtwtIRAMZq3TjXBDzm3X
AybgCsnNQ5acraHUCoWoRd73ovVTKdk79NrxgqpYjtBjBOGQozLh/FtyHyFedonB
keR8+y414pt4U2DDVUutp0KrSbjG2iY4bo7xC0QAhdvFSXAdnj6AZCdGJ+M8oxY6
35AXfa+0NHdxKcCTwhPm5xrYcd5OGDNNPXShPFYJKa5pGeP/4gnKbEKF6pA5h0zZ
MLKcImcqCXkgkQlb5o7IT1eLr8GeXe6cdISgf492YFCxC2/vUU+27ORIMA42pPL4
1qasB+Cz2P1Z2VSbI4lliyjjuXO502cFH/+wL9B8qq0UY32crnBmuK0I62jLPHBm
VQnQfynoCVB8A83DMPMWJj6pzv4+oLYLm8lgo48FA2yMZrc4K2naRYl1sBicRsaC
5w25FbfeiM+CuG96dnQ1RdbOzlCy/YRpYsTXY3AjMPinNf8eKN96Z9p3NOGfgvNs
Zy1HuvI/u7xi4G/7Mx0Yv3IedQ6tOpQ5f+2qVDJQOmmXreCVNbqhbOSOQk5XtKpl
4nZ9AHlcZoeot58hbnRcEtRTyI5a4t9EpVUp29df9kV1rE2w+LT5GG+GA1B8EsKO
BkEvir1nWocUD+pjdUmbgRgxMJ88t19vhlv649grjH7OkZ+oelri39ZC6uXXt8P7
lYl1CnD2mvQMdMyjFZEvq50SgehBFomTtDzr6GYr8p7RPqeDhozl+6rHtouewYcM
y+0qLGb4dseTzVtRNoVhB2GBIwL5E7aO0R7QAMLfMrT/oWqnFOh784fkHlWrK2co
e+GjhanW0w5X4ljJonobTcEaa9fuigXAs/DflYSmBhRou6KjEo1yNpcXw3Bfz/JU
7JaZn/+sF/widY3c8klSfUWWFbRSqYHO949x2LmY+bg1d7bV+xlq5M5+V1Ohl1bP
vgTr365Sg24qdxJ6MUhMgMbsyN+s7Gc4V/MkE2ymxbYaidNDkOppn3MSfrjhohBN
20MsktnN8GjFIKdMehlyVzaG8JYXtJ9FGu47TMQchs+hgnPwH7jfJToxytsxeS9j
tPwqhQhaU1+P00MSwi9jIGN12ECwlirf0QA2J7w0MiZdmw5YqXxj3ikT5zjiARRl
PE/X7J/MArxzTJ69ML/X398gnttwJk0/bdAmCpXnhHKM1GcBWl2LOWmqdpTiHIcB
ybC26JY8vOxN7+pIRUbdSIME4rLY78SVXjqqdncLQd54aSpAZGagIDPf2e2Z8EHN
V09niceb7njhYWN3ZjRJnjXEN9wuTfuFBMUc5Mvcf1RBUekO9R95xdo5NZWx6QAJ
mvZd6auSpxUZTHqAJx01bBcYL6G0UIh+UA+Bl3kbJENK1tE5mGQD1KtC0szfINbz
nhxAZJ2a4Cu1YTrNMwBrPn/AWBRCRkUs/HJgA8ZvT3vUCfH9C5V4T2P95peeVsl9
7FfpnPTb2ueNDLAeVvgBr2p5SZEHmYf506ttAVgd/jG2QxZgw4cRKjhxUd7EJt1O
tlwcHFromfPeq/1PhOte5us8Y6nGQ2KjnurSioBTAjBUQbrQJexSrAAPr5ZSgpVD
o/pMur9tZ86LCsxKVwje+ujdg34a8lXDTP30zD9Dp7SdqaW9BeWdODlrjTl7A/rS
E1Vg8hXXlCenA6jhdO31Lq/BxrDViD/l54It6MIa6FK2Soz0IOzCZCOpkT9S9AYK
jT/QCxTK9380Jjy0FN+zw0J7zpQ7ugmLsW4lBb6PPw8xari+D5at5SesSa5iGKSo
1kCPTdSU9eVivdewh7lUCThkSVpwA6Q0MLZaMOtRlfPv+N0rjppZB8ToxlwYvbxT
i+tPHZM2au3PQ9ZTDupHB8TP6suNZkbVa6oPtgMLgIUpD04a2EzAPMX3icYMqapY
JBj06eK1kd/A+50GcIRQchQ5rlRd1ODieau1FG9FG1Eo6A9VOTPhBGS1AcECegL+
r7K7yb14D4GK6GY9ZPtpV9gA75VmCd1VExv32mlDLedP3H8In+s5t3Hh1J2RAq+d
YnuQfIBVuvXB6dT04rnQoiCh0Hr7y2/go4izAXdZ1p0szAJzYFZvZocES/O5K8fr
p6fZa8tKqYRMCCgPIKLY5p5yfRgvQhyl3gAyh3cey0kQ72UWY7QbNP1w27JIDMXG
yskCJ/df7dv0MpGbFiFsqzm89G2PtjMMwqrrpEr1jSaBfCbMbPq1GLZTf58X29IQ
kzHamaWfXSdGmhOmN6bKqY1Sjvd1763veP02Zydcq5jdAsYVHIDhSi1Tcgm1Z0pM
no8eTGqdnR1r1tRV8YmNmGNncgZzhXtHYS8goH0BH/UaThStc9zDOJbai+4LOBJ/
89362kU/Emd0ZiK1ZluG+Y6vMr3s+JkbIvY80EhJEKzUqUkAyH0nHE0ZHTxg2Bkx
i6Eb4HOF2+cdb9pBzu32/AFa49kFtKi252SAjkShDHMkgRQiXGkbgBynfKk10kud
vONa+aZBu3iCUSOAretNQwA334GN/ewtw3V+W3GnS+o6oZiXlRElSjHgu/0F5gJa
phItlOnM/E/axOO0qctK4Roo5lPHANyCwr9vkf5uNKeK3hObINIss3Mmt2cuiFef
UqxfAQ6P0SJ/gTIkRl1FFLjRtXXAqeFPzapGR6LbDSiPMldGhrp9D+HbXD8O1yB/
WQLlqbFXPDAXWPcJvcvWLOSMdh4/rcqQPndN0USpVQR53QXxBiRJ8UpmZenLcl/u
h37x5v7WG7UpBffwWUWSHDGjrmUYhMhslw9JgJfrJvanbd2fYhWikG06FECpFg+W
G/o03z5ni11Uzl+b/zGxDGMSTNjcu/n7lIi/Eqy9LpWOc4m/+W/xKqcuJpFLDEzy
+OLfR32OEP03dZkubqT40CBZtJdDkh9fFLX+zst3EgkWQwZ2CQX6zDaEeHwC2Pi7
kdQG9ZW2CYwHNy1oGROE3Rv7YAFs29Rzuxlqg1YI3+V3BF4/hBYaSpmJN3ezMvkY
0t1B7KNa8wbfnSLrp/ZTkXtMA8qvnTHtusr6278gJ5+tQIxjitKj/fvcevLAkhLk
V9i8/f3EUW1djlTONqTdD0gxj0GXRk1OESQWKlH6fFOP9lEcDVea+UEn1FiCgYR1
oSnHQzNqaZQx+UMz42T7FKVHyxrK0cBpvs47/QTxm5rrCtm5BA4exzWjVBstpJCg
bIvRDOXM8qDZdKo3wzIewniqgzIXz79iMaq4brsyrhXgWwCJv97NYCBc11cMvP3h
9VUiyAVm55UBntRtFu/4EOOtWKKjb85uevn+AexrP2HfXyFeny27lk1MsTQbajSW
k6icGPTSVQ3Oc7WH7+j4uMVNg0VowPpjQuMSIiIJztWhvE60DJUC5nooZ8fmohd2
XDNI93MRLFgih66p793PeaLmyZ4EEUz6JZjLCpLanfBXUFHgdRz7+8tO0/B1bzWr
DzMnNLN+Q7+gAmgxOVBclvByGy8ri7Vco5sJbzptAus0gmwvLbbf6A739YRgdN/z
gNhRwMkHNopw29K/qiZInaQ2S7AP9jyDhGSjmKOfwJvo+qhp5DtRhD23NRJOSuRa
7gxoVFvwjScVyd44Pp9bj3xETzLzk9oBm5LMkLPk4Sn9GcPLo2wtbgK9jLxBubyD
0E6AAkrfLk6oKcLbNZMfAEth3Xq5sJd5GYsH5ghi13mmRtJRucxBvoaQQ+d9J/CG
S0ViUnQFVGXDLvMR8GmU1N2wL1yiGTJQ74n0r+zhJUGVEYRXdx69S+eFUnSgCgQx
99iokEg2WQ9NdnzOJBR08bXklbT58zlV3RsiYaKZvsOKGQICY/uJaQf2lk1gRvze
eXLwiBagkaTe9F8yR8bxT195XADdw6GuExeSOBJbfyghPw9qbC8/QmHVH+yBQM/T
xR0Bm/BOBmtrKL8i20qo5IySs18cqFFcMEB7FgGmSXEzyLRgNYLz6p8Cubi9lH+i
HMqa6C1SawsM6TPdAwgbytgxEwOXaQWvUUAfZxV36i66TnycPrMZkk+ZoZWfPVTG
3k8NcckapnE7+q5I833irXuBsg9IJAGTAfwIu1S92IcQ1qt42s9xUdSf/lHQwrKr
4bR8zs2tO/prEDpS1Jyerzji63iRFXOd9/R7l7niYNcmJOYB+jf5Q9mbRBxGoT/a
u5K3yoyr0Eyse4IBSojkphOQXyGYKqyNjDZCciQlAJh1658lfGncK0/v04+enVpf
t7QRXYPxKR/qCkuse3+RORp7SHGu2D9rQXVa4+2TJCormuggTkoENjweynw3zdQE
7QbSnjwfybP3ylcRxjRF9wvhewJnZR97gf2851BDUIRoQRpV2JTTZxLUg0L7KOYs
IdcmnP6nwkPW1qN4ZmPCZioCnE0tScVXWG+4Z/Rgy3cfpG3J5kvwl2alftCcIUBU
eF8OlPtb8aMRM+fB2wU217nnGVWF10kfTcJP1+cy48PiP8bcJr/iUmceLEpJS+qw
T2le29I7/xhrbEL1Qd8L9LIh0KzZtfntKhplVDLTetaUWZBNfJVlttWdJ1C96AYf
qU8FTGEorvTzo6s52BG1xvmb3sSKdZ+OeTFsl7pttp4DMQJFpHNvB2JdLn/Y1Xq6
P3SijbxKjyE+8beov6z7NQH/aKrGOFceW4N1Dza1rgh1YRO/g9eh4C9t80m0IP6q
A+XP3IDIe42zWlfxFH0Sy1wAmvu7MucIyt5wYQvbISVYVX4HrZfi4JZOCk5PR8xl
SBQE+iGLlutSA+oL8pJpuR2oH6m5UjEFoBCqBG6MmpZT7T9eUdyPf/4UY8ncY/L9
hLgTHSsYeZo2ICZFH8/agV/5eMuwFdxvgOFwUewcfMDmoj2J/VQfPKaB5Dpb0UVS
IRXZ1y0X98iIRM+RBUujkLjtfdMEz7peffNDjGXtIcSS6UW+q4dJNqIh42iBgH5u
8Rv5bMYInjQwQMXS2agYPudUS7uUJPfzka1CiHNw3zouSienIc6jvViE+84EuRso
2qgW2bjliRaqov2vY230si4l2Pk+kDAqOaiwoeVhZZUNsQm70yYOfaN7ExP99zQj
R+58hlOcBnNpaU6KkNSHLgFo6r+bh56IgJh9p5GtQFuCIqeQd2gnT8WU1PSN62Ty
XUgNYwd6+oQrIJG3x8FKBE/DszrTThcnU0YzI9drfb3M1YAIWq7eq+bMTEQ8EiPX
I6qIXxYIPcNl5T6lxci0+3ur9Mraxf4xKde6fX77/F2xbRC6MVAbIFiLyBxfiyfy
DiVBQSIyqaXjfxZZzORXhqUD2bUDJ5jLXiXuLqRlEpHwFEgzAF3OS8PVvAKyKCc7
1SwDmMoya87qhevidbYiCJj6mDquHLwQuVhF9goo1ImFOoXD2A8dc7Fz6ntkfDXq
9gIDlOp9UU9oIfKW80coUjOJ01MHf0h39awBMc9N9DG+zFzUQgWw/4+U/2wMOpHM
K0HBLloqYonbB/+GNdWwUoVwgwmq92RYEFL0F+TObbn5IND0PCsbmLtxbac7dswT
mNDcSU31ZIEEBxU9RheSQ+f09LBlRVfzj0wcwvx3xKcaR1s+WuUErDQEGIYuh0MI
7Je+c9EZM5B+EOdMnjasVI8tt4qPhRUn9iIsby4iCGXxt72zVttm88TVBA3kTSVp
DsD6CURmKL9MqgPGw0ZkT1nTSm1C0P4nnjeqnDHCqYbphh0GJGj5EjkBRvUOa10e
aTvFOITMP4PrDb4tN/JHOZNxNedNFsIP9Zo936Eg68tz8SLmT1nEWq30moWxrqpg
g6BjeZ5EISa889xADchFAh6t34FuKYfqdhTa/KYIzUlwL+7IJntt+yiKF/x7JsGD
WsEtNInHf2+ZRRFNDzFzwY/VnokkaKqE0GLIApzlaagxLbBipyizMRSpJvQ5Y9VC
LF6tOAuc66XvXhVQDZgrcMCcz3mnyD6Xnbi97yTgqK479po0zM8PA4k5Or8izoxn
gpYSOpiCoYD0rQf+l0PUNK31mKgJ7XKnAhLCC2L4Rq3ZUgAm8X0VRdve0LKJ9pWs
FSx58Skz4PGJgNpGQkUrKk2gBM54WPzaDQ7HzWR0K1ECelDmo1jBFEvPGOdX3cuJ
oIbjdWMW+RSSK8S2UkiF/v3dLdna3Oa4iwult2JLkOTVCQRWyso6Y8N1ITeT9oN2
DZAiiGsF5oXzMJ/xyA61WwvVplZNrOQAUO5RAqBoYQjodIyp+i7amiKcxgORZZl+
/8VV+eEOEc1hexKo+X5TLzoyiRDK0jWSw/3YK5vIhnPE17Hh5PPQm39qBIMKKWMv
wVKgjlFD/rEGRbRbF24wFFbjaTRWG17jatbVCYg2o2+mMOvIPXxKUeDTqerHWbPy
C4XrccBihfZKlEiocWahlkbOKOip2U88wm9DycUR3qBg2vTD30KY1FilNmeMF8zf
WtJOqAACu6Fiu39hR32DZjpY6p7/0B0MfLNEld0oBGqb1eFo+qOiBfXUdCRICdVm
nhwmvCjnktA9mZwfrNwlp+RsR3INWhyfsd5v5boF/J249j/BliNsg07y+tEhBGaW
WGei3WCGXp4RKwK1vgSHhYDtx0QOfHQbvckHiswywdlZj/kQkvv3x2YewXFB12zP
zs6Yb05ELhAj250CHcoROEpo9rR8JTmMbmxltm4LMHuPAmW6r+fqPkxTk17EYpfc
o5lTZsRpaEh+120H6KJWAADWbUrpkhOPpSXPsMVO9xP9qPMQb8/4zXh63x/P15OK
GJmXSojAsIQ5iZqpyn4vqKsfABVVU3lpt2lluH4md7tEFO6/T8rTAZ5I7cuUSlzj
pb0na5HpLeC+ccyqINPYWS0js9CM5NzcagqI2NKD14K0ye9YCWSdYd0EbhlURoCj
Mc/mQiT0CBINnfendZBZcEYoGQWLVXQ7Kn7HhCRf9Drl/KGaKd9J7j4VYH9A7372
fIUJ23VaucJvfvzRjOcg+tXZqdMkD4qf4NWoGom3EZIAtW0UIROgbQKH0RdnTz0h
H2ep7YhZUHHa3K31S+e0Q9Tkf4Io8131jBYWrLPwabmVuZnwMhFHb4kN7GM03fyH
gYkviy7hWcSlDecIBCafcXX0LbrPNRxFuwaPV92oG1jF+sboEgn8ePJ4NYnjEyy2
F+MIRFOeGjkorMFpCetLSv/YBUo9V9+8Y/0jnyh0Txr6jT4tKpH1ot6RyGOsQ146
5HS2IKko4XxDtcfhQF7WdrKnlMEb3uaLtQaeOae+8x43a6XUqvat3MPlVk9tdSK5
UKphu/06XWUIAMOXGkbOptrw2nQczMxkVak+oaI1XEy8DzSI3Reoq28ZOrhvku6k
ch5VuXNFysgpEGBdNu/SSvJY0f17fA2yb1sIVTSiZE604YQFWXjOSkXe9/jXO25g
ABtb/p/sajxLpk9OzH//72JFC64gyPoj9+7FaB4vbQwR86uSM3qpD1jhYiWM7hgG
mSaCjEfkKkiIgRM3NRKIAYkTgCRohQf6TGg4oPCKiAXT5W0cHoshDcFzNp0B6ELp
OY1uwnB2C9xCwjRDK1LwG++IKzHrpNZDBmCJB54f6xPrtRboWIRyPjSwuoajLjEw
WTa+Cw9MueFKIUALMy7SuQX6gOkLzgyGmAn4QS6A4sZC2Sji9avDTYYxSrXbyAfr
0MM/SbU/H1FHZUbKWlm6dp8EQBsRs5CV9T/DB6Pi7cevMOaVkGL/VUxKpx6LwLtw
jyi7s0THIYP/i3XWeJB0jZzHSREYHIl3KzzBBhZ2QaeDmk2V4GZIBZzg/tWU195k
HTiBsWahAuTLIYH6wqP+7+oeRpJISIdgFXWgReD8GZt4Zr80WCH1SJtkzVVjeKjz
98YVJeEQFWSTMA2/pdyZTzKPNLbs1S8slds3Vadh9xOMvUrtJY2T8Sso8J/lZZ5J
WzOVI96QpZ9VvUbzcoEwi4NHWyoKfUB/is1EpUSmSGHmoanNQVkCQa2EwJJ3Wcjq
aBcNpvgDwmWThARiNS8kBOoeNHJ/YP4K6v/qjVZ8WQShesuzPID8hZkkm9vATScl
7DSuu0bYcJ2/kMUs9yvDqpaoNoiXaNKV4Gk9+BJHYvuqTyjJy4ZWBZ0kI4siihf/
IqyV81Hjr5V08duHw10J94+fQjrR7QJJlnFLtRRRE0EaFnzILn4U2PoTU+75nqFA
+Ig2Tqzv4JnDRwmREAmZh4f7ts5vdNpUiwJvC5Rw9z7Sp6Xfzsn+O0wJa7CSZ6mo
LTbe/8ClFOXKbVi1LrfXFoZByTpmfosMM/v0j2xwNEKFV61WWk5MW+Mcuxhm9yQC
mpGnUE+WME5/8JB4iZ4t141Hpj45DjijSj8y22E3GN2tUbN4GGx5TnjeX1IJ6ruW
dp7mjjjZXIeyBRsgNBcHXILe/mrOXG9KcsKfOCDB7BN0C+DhGEyuY8e+icGFskcw
z/muiZmhl+NIt66mOgEgcf7vPgIMfomd2QLeG+ifu6b0oMkfuuLCTjKTz7ZbhvO5
r0Hm9EHAjCSmmE6Yo9mAswxvnhLgSKBvCivoOos2cLg/pwt4tyR/eZf0Dtjg6JYV
YTmAO3YvtP7Qs7SqzJMPmAGqwF8nsFG2rPuB3AyW7n8fZ+hsyLxsHU+dPFw7ociU
Er907wW0urRflAfv5akA0pqeQpV7dSuyGqCMPYXYLFhgMuuhL4z5JDDq2E0EGd+d
Myt7kEj45f7/+Gweg6znUCMEBs3sCi+e/3ha9V+IXjhAslWeWenXzpSG2kuFGyD5
DPAPi/zormfgdCPXjPk2bLGxo0dHamcgUXV0eLXvCfEdtPRWMjkB0JgUSXXTZ2Xg
KTuT24Xi8OLL/sTkHZx6QU1aVfCjpKLUs0cLjSa6yXtztqbrOHe6W4OryJ7n0eBZ
gbxHWmZK+59P8bbOmHCvl7wmmAiYh2bKvML0pM+4BlOG24+fJNzNE/I/HC5dFf7Q
gReQD+gSJrHr7Qoh7ffSbvRiYYsJBtBrkDZM5TSXvjc89Ulf5c1qfj3G4JT8ATpH
cI6FVOduKsMTtvZgAukzAdwY8meHtXdYhZIN6nPj5ongffi7BdkX1kIrvB7CRFlw
OXaeptx+u+W2wdpXGNJvhygXdhCVILoarexVS5tyhp2YhVxsZIGI18uM6V78d+fm
Q7CbtsFk20Ze9jXDpk1CyoVH4vse8Xn8jqkL0vU01mHp3bJ+MIjZzgnrx5w5f2jK
TKDYLsZwURN/iNLpi9meNckRLCioRWvBMCIj2hgjA9wY8jXDe2oyb/rBXFeHHAwI
sjgNcMdqmA7qwuhLWV7krloubFAlFfWsIzB7BigKS7PtnjvdDXi5RERptEuqQNtu
cHZ/c8dY16vtiU79NkrEByJ2XE4K7lagOPQvzNNT4VYd+k3oRVBh8caKmRdtZhDI
8y82/PJZx55IxEEeiO24+fiCP2QCJHh5IyB07ydRpSkSMc/sWErYZe8EjxqDD3q1
ZodktZvhYHa6w+CxOG4ohScxcvzQaWA4/P/6niUct2YaLV0WRdRD6dZLSirnLBIH
Lx7Zzu8HpPElddtTnTo4J8QS2VZ+rXOjFOOLKlC290QMUqjN6+d5p2MQsEIqkPa5
e56VHupU+WNRllMl6R3oynfGd6v7dqz5NxLSmtV/wl2ZV+RC0gcPhoz7kSmDoqFy
1QuMgBFa3HyGRK3BiisU8Bh9e2pHvC7/goC0YMApTGe+gXqL51JHcSQdJ6RvrIve
VDMaTCSZyUkuzxpvknTNnBJUz40y4EHBOEtUvXdtIURynw48ByifACjYajktE5cU
M36/H1IMpcDD7zfZ6VJi1lt6bycFYoHUdqzmdNTb6T1B65AQ3kq6MJHAElSCmyoX
4KfaYmTL5GlE2yVj7rAFWu5naLpXIPoilcztUqRJDrqyh9JjOSXgyFJc7BdcxnxU
jt7UPx0N5LBJzbbdU8aE3w5oByF1g+6hL1XCDcG8De8Eqeio70+SQ352W7rofE0k
IxbP9tX/S3DMhqQyz/vpFPj/Q9TIcUHmGTHkR+JeDKab2TCUqmS1d8LfzwCThXCM
fH9qJxDHl/mk5b7a3E8sk+qCyV4GHEFTKJwK/lA2OaBtec7FN/VdokhSfw9IfaxT
sL4cqq9nHQt69ITbCjPOeOhaKVF2x6A73XZZHznTs2GJkxoTjIO4t+olEzsZhIo8
Qh3rcWziK6/f3XLfKGxRUgDtwne7UYE0My2vj8N6DiWqCS6c3AWQYQL5ubPndZpl
I7SsI8ifA5egd+H5ERxhdkA2Qc2FdZRnrVZi3TGuy85FXEtYFcCmhDq1AtaJN0Te
4FFSRwfHuYOr56TV+3le31/c2KDxyXgSskP5ou9ZKnh95lHPwiNB47DzXbQAofj7
mNmXe9w7UVXU8tGPo9u76N5vUmZT+ey1xwEsAfamevz7W+QmshY+0tsm3T34P24z
kAY5rmWTNxSd0wwO9hZgJPgY60Jf1ujvy6+Nq1LaoPYvHeBPqpQG39ARM6LOwCeP
TnYVroPgrilCT178Q7hTHiZGFNlx+kkBB8xId8pI5405zsqxqNnEDsAwBHLn/kxu
5JG2Sga2UDFCrkjZXOLZjddwYf073sHBCXCBC2zUfBDwYMsAqj0Lt2uzS81iiDxb
95i6PLv07OcfLrW+4oyGF1GLgnrTPBHgDYNmUyzSpw/ZMKCFydrl2mpuucVXvqq3
Y9X3xMjXlH/mwOG5t8S4ODt+ZBvgn2qjG6wwgO/6i3ZrarUIQUYGRMDCiE8PiyH7
yRfZmL3NdUvwNU4cJECud00M3mWA2fiZM+Y2IDlZOGO6GsjWVvDnvMJh5H5D17xQ
25C9QenamiOUhX++fkzYDuvNl1qiPNw9WtfOD3y1uz47A15uWywqhsW6CparxObk
G4KmCZm8oiKullfScam2sXHmmoievuhGdhe+2Jka7wDe10EdP4UkFCSDVegaQZhL
22pe9ZzgOsbaCYJFQC2mAYihAPbhyaDwH3UtH6lIYXnK3d/S2mKc5ViYVx7DgU99
b33po1sDjFazYcq5YWEeFB4/e4FLOgNGa6DKo2y/BCrdocT13BqUonOL7dPHeCoF
Ok0n665fhlObXLsAf+NPEju5CruBRcFnQNjJKsn18f4BgaxSYKSICEgK5Ep+A/wQ
HMPTSwYe/RjdBOklsZ26Nr2Aqe40vUY92ZcN3fKW34m04YtjHdPzBOOE7UdnlidG
ndeRtSHtutvAX8mdcrxqXJOFTZg2rep8qSvr513Fc0dN2WhVkMBg8kVc6ax/NYw6
EYHp5VoZh8Xi5h6ucb20d2Bj36qLsZfP3fwhXD7wfrXjD92cXweh9L5cDjR6qpO3
AtlgDThI6bCx5psgDyuBNgvPvJz3Z1rkSAxRRrt6+GtIuUuoh/GKaZl5YYqxsyIr
LA2k2yFyKk4CAH2hvjEuPmBniV/yoMrJgec1C6u9vUt6PfpGD4jKYN08FSU4/fox
X2uaVdeKpXHN0T/2AQYSbv6ZKz14b6LArtoQkTcSmAWkhpArPg7XUYbVu/WqzRhN
9B8OcoQcY/JAoK+ZW9oIUUWtBYIO2xER5cPBwaAllKKiW9yMYayg1pcsiw4jaknH
5JJ8Z5jITNP29MPd1MZ7iyY5pXLqVKFg9sFS4m/DzkHRQYVZgkKjJuWlFr65mIIS
cQRwPB8yb2aCjn+RIU+d3vvy+oomi7A8EHbjriifJc63+Bs8APFS+WUW8WECgX1R
KCTV0JLROxmhhEB++kpT9E7p6m/4Yp683y3F9mtRgeafP39cIPBTbh7mcHtjgyLJ
llvbbyLbftY8zTC4tpSidY7dUcIbephAREy/OwE1tHA1ciPKdIizHC7//T7A9+x7
uI6bd/ZDBYw9xTJZ0pxdi3+3RT3OSc/navz1N9hF9fEOXLYlHXR+j3X/wKBf8zkc
mXJ/csgsxcQ9MCDTj1qNFhBTvcTznoMen98PwC7vzAiAcx9facGxrAVFI/RF/M0e
+PIr8sJY5jiPLmZwF4zcYYdcXL7XxHPrBG7vaRHDIe3NFUcUWa20jd0w+SI41s/F
c6FAISiGn0kPUd+gDL4GPJduT5++piM3eobZVX7/oFMeHj+17x3zIGaRBl7jIj46
b3GfclArr+7r4AQDmZe6KEfLR/gpD91P6HyEGdBmK5Nz+u27jHVF4wVzGR+37KY7
Lh5l6i4nQy+5XkqfUMrq2A/D7BD9c8FkqAx0lEtklGc0n9QrYEcMLXIzDx5KucaN
fU3IiorMk/jts4W5v/ECEKO6e5wg8dWLqEs+t5bPZQfeScYzg3o4STxzOI3RQTN5
HFatca+ujt+85JmG8UqpZQwEQyGAEYHiSif6rfjJDJHZV6jxe0cHt0ereY+IwFBT
FZNBEXFqYRCaERK7xZoKFlk7UIOY/JZx7LDc3bEsWWR5otNJqmGrrLliaBPmZgW+
S98ZpQ5JzDKJ7DK/MWNtCl1qicCHznYFHZU7eCVfhwq4LMR8CS9+K4edi7iT6QL4
Ghd6GxV9NvEPHOos+oXPBhu36MmUqWfOTt9qTH8EXotpLWS7MxuoPL52Q2fDyJop
cX6ENaDqjgGKfUwY+cb5URGnF5E3CEidPItKzn67JheBw38abNJhvnaLB7OYm8Cq
inPrW2uEwna4uVYVpnINYjZef9uOX+wAjtQBRAtHQUkgKwtAOBoLEEHlxCteodg3
3nkNfpap5sw29pwGhHQ0QD1khRNGcYW4q3Iu4H2Ns7OlkXlLqcv9RPhMdQllWKzc
UtEZfgNMFQfsmkbJx9Bcq9MgApeS42ReCaqx7DFJtcu4szqVkn/8ODIQgdyRqHEs
GYCiNG8apL791t+MB6GMIUQQh22QugEquZT6G6mrjPPhs6qckKhYI7/AdUXdvct9
0fHIGgbMt82utyAY2KfReXgmqueWPsJhM68zPohKtE/JBYB0hy+ZGHzKBRwn2Gmf
WU9j76WAAlqnginYwovGnaMI9W5M232tlyGMy8ZV7vHFGWXsp3tvK3owsVbA6ybU
4PCKwFkeQh45wS1AUgkwk5T8Y3kYL+CRngWEh09q5FgwCDhGy+9gKKVuSBJEXdHH
yTXw2jT1+4O3HPU6tWu54T/Boxn4vTpdnbFSDpm9fBnQxgmsdWrjDpCxUYIQxIoY
dl/pq+Kbb2WDBEXCwngJYymBe3LpRskFiC3xOTJkNSEFg8Y9CzXjIa5GrtVUjPTU
buNewHEpgVjHc94KDlEX1tPnhZtXX5FLh6DIGVArcSpZXLHRT5/XR0NhowCcsRJ8
2ZQVQumujlsPJfVZahXznBrxgWYI5wnxoa5XmXBpyND8Ts3Kf0mpk1hhBfHnoWol
NDN2MerYUIuyFG66mX0eDDmdy+Qfdv18Bgr+f+rIrTSvvrOXqsLunleOKLO98L4X
f4pSWosEzGxOBlN6UreSO5Y1nKpsX7s5kKt0E6PIcwdJ6HdZSJJKrJN82xdwGjFi
tomCgdB33Cw1PjvgPP4T0uVZIFity4q1Qemnd8/iuHuuNnTp+j7poZKQNd7ei0iG
H9s5bB0nJMXZK4IJW189Ru3D8vgXRb6yhOhoXbhJMqS/j+Yy/h74UdFLw2JWigif
1mo+C3UtuiJ4WeqMZa5U7/x1nd14HQNXCFwTM/5NYkd2/SpgE25/K4q3pOKDAmtL
RKrm1+FO2Xh4zm6xR+OwNv9d/p3AjsQS6ElmdwvJER7R4lHRM2Z+eKcGw+QDWBeo
0JricgxcPx+xsmi6xzuPb36tYw9fVm6ry/acuV0BeQVFJES6w/N7UNBpFBvDUk7D
ip7rvIcslXmCVd01cSk/54pEEIxmYPJXKxmMT51IYx7CiHK/3DpRt48C/old8DEs
6JwvcRUrbnoQ7u7RqRX2VQQo+pWEwrn20hXW8U9uo1hdxlHm3JhAFClYvDs8Iasr
WdviK3beySZxCJfLezRYo/tnvFujIYUTY4dsVN8o0fNetJFVfKumtq87P6yu6nOl
axFTXqtuQEPcUFBu/Q7anGaIlJ5MvV64DuMhd59YpEPq1gYOAocY8PyznCLyEVaJ
r39uPZLNIC894cv8942p9UDq+8rvO0PNmr5Qq/MLrUGTdR4y0AfE5ecxc+cVaBWj
Xj+AiapthubljH2/KIhqzPQul/SX+ggDjg4JVSddwopzRep+PLK/j6eyqUMpkdpJ
i98tqRDoGJMJhYE7w4EFZ/8HjWSm1NaYuWxXrAlU/I4tAzcQ0XFBaeTmtejKNiq8
OnIbMDbczAV0j7ySq2CpcHUwp2IohhzMVhwF/BQlHUn1tmxvQrlGyKjZHNl4AepW
VKyxIU656zn79IvRKfOY1SfTQ2NTOZsdF7XiwGh0JJWameJwytyr6cq8AdMj6lTp
k4Wtj559mpsZ+DYFTCCcFG9idHH74OMg7FHR2O1I1yDe4QaoZot8jTl0EIFAVSIT
ztDBtb4hIyRq4PIZxR1rB1vQ5KF69BWYo2ykmvovA24M8gGcWigWYTqTqTUYIoHu
IGXStdaZk1vW0Q/tGDYexGIhbr5HASfAQOt/4XIHXJRvGW8o1u738ElrFlkHPLVD
J6dfecSuEJC+96G0b4ZW48Wu4vcGSt3RUTu70S+F+vjNfLwlV6j8JRkqKaXlZPuL
3xpadbpLW51KqOEnzO6rqE3CIO8XIxK6Qdu6H+G0aA6Hg3TNy2GmJXc2lYeaFOcl
oTYHgF/DCxj3oR9i715rMuM5/UbrrZZNbvgUlg088onliFHw2g/f4wBBcGhDaC/L
TNFWrgOPiNgKMXO0aLHXzBWY5KbVuT56wRSZ4poXnONdGxFi1j4vak9Pqr8iFtcw
NFQJy2U3LE9m9v2ZHvQA5oAUCAEo28XFpc6/St03C13ZFdVBo7AA3AuqDPxnCJ7g
hgJWhCHTBoXrMvtNkM8sl5DRwXmHkfNQhsED05z5lLBM0D4UgisxEEL9I9oy+8KV
QW4sj/IH2EoK7lFIyIAtVGpwLyU4jmWKeZ3N84JTc+M6WZmWTxAsi5OJn9cnhPFQ
kyZIiLK7MBf87u13TbwlHM9cXqdWE/MD+AD3ciUnZlsjfVkDINL0/KBspyVbVRsI
+LkmSrDnpPaCJo8Lo4KWRS9yZuA8mwo4wkgHHr3IrMZt2gZTUo7W5PzJT+D9HBdp
/pWADHjx4EpQkJ9SiP6HHic+QE25J7r8wFOd5b8EjGSF8zFYeLDYYODLE3CNRVrl
AThC3QMKa7LpGPZOT21sSrYEfFW2OxRhu6DF+Aa6tmz25reLb83cIJZKZh16gd5P
NgUWqyne6b8gVPpUe9E7AkdWV/88glSx+siF8d65OeAsIqu9rnAmT1NZJfZWFoie
MqhIyxw+yy70L0ycM6C5XnOuW5JA6qvHkhS3dax44Y3j0Oty9VDrRAxAS9ZgBuBP
v0F05nmo01TfuzkCenBC7q8BXkPwu4W456tikqq9TdBHxD9yQ4le93p5jjazqnGe
hJUsfEhBHlWuj0BdrumS0hJIN/9dZt3/Ys6TYWA4esGGwhwoCya7lySJXpv7Iea5
RmUppFlU9rptTeSoZYDS2O2wrDmCN0y9zu0OrE38rheun1XyLssSrdIL1h2UsQly
onBZqJFGcMNO7/Mca3ncqaPqBDtVuiBnTJUWgQMf/ZYFkGsHQnx/vk3rLvbbZumE
gLTvGrno78WvrKsgO7YEzkUfsjwuA/dg7yV1A/AvrC9948D9XJ/0SR7vq4ubg4UA
PkosJbaZz4Xw+LYz0AYbErixvOMDWfp6Gv6qrOJHx6zx9StjnkGMqecC2EWX48eY
G39NaiDNV4G78X4JE0pDK2JMLYm0ICAfp5wlzJZa8RgXFx5cqetUrdfhhcpZWiUS
xX/VbMrNvYzlkAS7S/3RcULbmIKdfgo49oF+z2ZSrxhUQBJPJj8HZmzotXbfQnlN
/FP3jNZJwcfrx8eITsn3PVN05rS9k0UiztiM2MB8+u/kc+u81RdwguLWWy3TYbxg
JKrsnGFu9nDteLcwHJj0elytx93STFyRa4Lu8KrCsH6HWs5aj9uPC5IhA5W8XMfg
ADQIUhbn2+fgnk1SjImYePqS62qaOIP1df4ibpxjpzOb/+JVjx6jG8f/JSo92inG
tQC1h4u+CUegd1OwuHkRsPUiWECdk+hIddYkTzjPA3Vcqr0V6B+JMjXO4o9Ze1xg
KR3elX3ueUH07GBmdRJq77EukS6/PvZwl2z39a6lLrin4J5WWO41w6nK/lyvM24n
OaRHeLsNWO3P6PnFO4aBftlR72+5z/Wf2qDyxwifVhV164KEsnfrdMgizsWoQZjM
lLhYZdPjJyELOxiw5yfDI/45hH5NfiCX8+6NwpHcbrrPi5FKSeIMS59QhVMTlmPo
hpyxcP8rBBRGe5GT7U8oLGkD3KzQaigahy5KNTUtDPiJ/o8bRXSj4BEATZakFint
2WHm582Wujv6++1r8gz8v9X4YT5tJmpHRXqI1wpedB+ILzhwSS1fE36zFj/Iso3a
UQn5voT1m01zQ4T3I6ym0GeQipySAuNxiK6hNsePgYR3S3bs3qlQrnCUT9Tthk5Z
VooypN4PFJN6QTCc16rNHkgk8K6bQAQUfVbsq3OyfeLqqHxBY1MRUcD8RG/CuqQL
U/IEoBCI2Efx2o2D8esG683w2P1Zj2XdH/MLCDIVhanDumiBFCZGX4SEAdVIzCiw
egYg/g8Iiw5TwDbLhnMvT2wth/iK3Othc4shQT4Cmv1KFaJrRxyVOV0f8K4FDASj
bogPQPSdWC+M98JDAsmA/8Id9A8VS9/tSNXbiClNPGer+ySIu+vrXWfGJss+0gvQ
575jG9sn88+i9oc+yP35PcGnd79ztoLG24a5K0KifNYUOE7Dxg988lj673PvsVQe
htVcpxkrNvTVAMOBJl9tgh1P+51xmUC4muB+Xbi4G8QcaI/KMffuW5UOQi4w+fUE
SC/MDw8BqBCnAaz0Da1wqeUtuE6dFUW1oJEMEnTNEOj9s7qkr7zUO89IITaIHYPI
1uZ8k3J1hPpjFyRBe4C2KfCV3P/vUhKcKJn0lzUu3kfR00htN4sHn0MQpTVcNunT
AWd0MJLqL/8Mt7Tzz5+hIiMlMbMdUm5qGSz8CZhzj8CSKD89AEhfQEddVoXe+FH0
nv0XBL2++mp1cGXh4ecDmVFcvmnw70a5PwgANqt47pcRlC2G1CAZYqTTQ1zCNHOJ
yLGo4WLUUeeG2nBBhOYyGd8Ta7W6ypGlY5MeRkHbCARkwUjmay71mKjPGq7QQpSv
Vz3UZ3khpgOaycb5fXzzs9icDZcCjn2zZ8PvoobavHnZvA6Hlbw2RuVOCZfZaah6
jrk3LJHZgdt41nfR60VvPJchBIvjBZImUzmN5Ko2NGw2X5ZQtKc4IRR1n0oJTAkp
XyffiajaT5hMZ0kVA2MYUR8qgPQT/jlWqaIzVQmg2UZ0AzWkaHm6M35aT6jnHPCs
66gXFQJXT1QCsk8mtxh1WL4iSr6/aqEvy0WTt+J0KFojcNHCCJ0+rmTBV3onBrK3
vlzqIr1S+lIRjEpwLzLZqT//M1cVkCIeLbKV+LrClIj5cg70wUJS7edxRWnUX98m
i+w8YSmXHf7d9srjH9ZJvdMzm2AB/GOvjngiBSotAkU8nTRp1CXxBoc/qvmALchp
Cph9rpQJxvIaBUaMzvp4hZQVQGDR38u+mo2vahdsLsAy1peY8vYaDAzoBDtys34n
nnXxwQDnQhvDW5ZiCbtxrCU42qItSRhCbqFB7RUrTtMwNACsRegZ5M2UKhOcfsxv
N3JZFeES8FvNGy3n9pWAIgaxu3VdWBWi3LdqN+isSQHbmcTfBIFlu6UZz2cyhxrX
vPU7gfzfGpYD3848NriX9PlLsC10BtRB1POvKkw+1iibGeWMT5A/8fg0bfNtqWTG
1nC41oUR7dQTgGg6r2N95m5sNkwoimgNeJzTIqeK/DO2efPfCk/8isQ2pffwcOTL
RR7DXU1Bx3ePJ0cWjh3Jwclc79Dbz310+e9oO4DBycajGRPZeKuw3V/MjcGIgF6G
Rip/FTO/Ll0zpr7NJB1IaGk7jLZfXmx+V1PBMkDsQGdvE6AmgJaZVIP47/jAf4ul
wfpamMOeJDz2sj98RT0uxrVl2gtIzbes4M6ecQMWWNE7XMiIfVVpVCyyrfwgkdWM
B6lzGRaRLuJnjJnQsXRCJScxyzGZrrBf7lVaRpeUU9SppgYhCKi1NFh11cTC8rbL
UCXzeTM0uDzBicSxOqGFN0AnLkyKqK0xm6bRdh71U6tT44Tf0rDMpz8LiLWBQzEA
RUmKX0E+NmeS5mN7ZYpO1UMQUmSeA8ZswDwMRsDtb5d/JHhTEzHiTjEoIC5dTVw+
FtE9L2l9JA7FW0U7J1p2AKBqRv/WbSovd3RgrCzs3l9KeSt10Z2/DzuMAmCcESRn
x6g01TXBWHU153QxUObl87Nto4BreU5X/qTnh7s5QzKT8/nYYqxp+yUxZFcQUSv0
2DyJv7xjNWgLeVTpSW+SFcGpwLDz0rUXErEI2HXGl9BfNK8Hpp3s8lrcj93ZusZK
h0QZxffoi8qcQHff5YzYlQD5F1iZr2sbdJ4YdaiGvzLIl9Hmy5iKfOsKTuaqBmA2
ahSj+fun5m0jtZ00cj3T3JeOIASEqTNvbIR5fvh4Lw4S/amyIfJBFZOPcKu1aOMd
8Bacv5jlshf6v+QNXpAKaTbF52JTUeizLF/YKy9WeQq2TrmdCDcsZQVYUim7bXnH
MaEQREz7aY5yGm63ijSZ+JKuxBUsj8Lua1nu5wyfm7NgFUouRFrBkyvulWpZkCc2
bIHg+TZ7AmPB/huH9TPAjiyPWRH5kCgxH9r1Hmty8DT4Ey7Im23qYOg981iWqOrj
d59se5OBBvrqRuTG+D4m/LMcLzuteZA+eTWqYLpbV66MH7wJ3DZTWKsCYgcFQ8iO
gymy1pI1Ct5VAzTiId9s6bBlcUGSXAlq2R8Hg8GDJGY5+0QzB4L0U3drXyIkyXLD
c/3LkmHVTdrXU2rNVfvRcA3GnDR9gqwvXnT2VFDzjpyNKZulDgZzl2OU3NRlQxgd
qQxSkFLabUUEEHtPVwE10QPVTQsZmcEHnZ8OEmmitSie7JFdUpn8xXyhMo2UJ3W4
c5nxI6hkNbqXBbvuLiklvZWlX/AV1ji8CDz7/hlvX3MYZ4H2229jRN4deWVlFud0
J64jTOpN+AgsU1NXMlGpX+WDmfPT6hYHmX37XSqZYhMxsmKQPcxXcvMm8B/7sH62
9qQbjg77uaCBHr9/UzSicVsL54y6sYeDDh9mDymSFOo8rVWiROpD8p+EY//LvaDl
N2sc5Y7MStvgYJToBIntFm/uQZOWkUu5dEsLgl8yTHj5PCe/X/oWJPdmyre+wlwx
E2x9gySW4Xmbx3ejoKDbHTNSIEgQjg7GxO1A4jAiOnDjpv6kcY7vrusFSs4ZsaZs
ePvZ763BlzsfDu4jq+WvEC5DaRTjLfwMQrm63Phw1bM1Uz5qxDTuD4/Jg3ACG4jR
mNasXAJ+El4MUZJFFSO3tHi9W7ALBj6t9MlDIFhh4Q8OLlTYtNcTo17Ttjf37l2b
/INQSx5VyrXtbrZvV3RvKkPxyUCPWMUEKwBqYNcSGLMrTg+Kh2I1U03LxkuPnV1U
v/zqPg3G1bgnR9R4HpOp6WzuAMwHYNuOhrVY2SbAPb0DRmTvwhbVwIwVPjKMyWTa
u+FIlt6+VXxvM2dciY7OM/lo7hF4esXx3AD9az4uwL5sKrHYLxgcEQzQ/MIKRdPX
pqrPMytNOIX5XcasjsqMf5t4qqvmnwFdqr4Ip70PTxdEF4diuaXT31XmXvuYrlM1
PtlJowvHJAmJ5eEKhcAnMWuM+wMRTekSlbZca9lih/49iDZTL3vunQNtRMiXBIvX
ebaDLvu9+Teg+67PHXOSktNUYa1jupUUrMk1XkaE9uta9CsSk0KC1Bl5c4PVQlZ+
tCfoDdEjRPfVb8sjTKsfrxp+vjmzqrZe+yYiSfa6PExEFfGe3C2qG0COEmPRejlS
31KgXWRk8Rln1nGDY4ICuDjrnJ9As3hAQ4upgBLEIfQZvMIf9fkKGIDYBu4WxopT
EAipOfoq6UAU0eE1/Yd48LXDjCG6RAVMlQmMixxh+wcAJglyMgmJFBYHOo3pnhBg
OIVqkepHe6jtjL/MUMUjwCBi0Ipex6LShH9miej7uigAIdYAXzRNWmewzhV1YZcM
3qjDvsdv2Q5deIgnXAjd95zLQOfgo8YKdio0z52Vun7QyBIWQ3PD94X5RlsNT+17
85LXLqmEj/l08MV7YDELNqnni3AiMY9TYazJlVnStdHdD5dwksaE0z4Gf2Eje0Zp
XEioLeTXD7THKiZZAlTa2Dvm+8/2d292KRQKe0q8fTEb4tNn4fu0paqD5QaFX6jw
ww8srzliBXfofdvR4NOfth2/bJBDHMJ9Y247XLGGMWQI/ujvX+L6d9TQqAfRwZ66
nh0rSvE+vkHR75aPmCtqdEsPgCKLQHcyRnFihE+P6BuJ43IwWPkTHMl3bI2YSL1a
TowrRvPw8GHHT8lQoQxDvxPUeyEQzH3ijDhiqd6IA5PGipHZ368N8+64lpZLwTBG
I5YXZ17mvK18Qwf4k7t46IhyZ7UeGkGgZka9acUaUCre+BQjXiIVfrEWj+o8BvjP
T9T4k0er6FBBLYMIl8yE4M6nus2E+xDc/I8fVHh+L9g4HqeAlaO1/augR+LL0kWd
HeM0kt52QUZ6I5YUoFyBvRjHyhk0TpBK7kx6p7baYy2FkH0sotq/hGHUsJtJ7Jdk
yEfRGKEYGscFCRNjnT3H1sC1YZ6tY/l6p2fmxFemIqaLZ7JzMnDEyrUmbacjH5Zl
/9PQBtoctKHtvoLMima/1pKIcxiM36+R6uWpZ8YqfUugRsDMzRxEhgqD7mUZ8mCQ
BsSD63YPW+Q/S4pe28dWBAbU7OiITA9kGVjlrU5FeNDUuA8nMkQyL7L/Tp2DE+FJ
Kl+vNSL3F7K+6OppUPysZYgv8z2yFdd/i+Fmzxm5s8+QNvhwdqLYi2BRrbmaH5LZ
OOz3QpyvweENTYRk55uzYj+9AeREkrrMa1NdnjSkRpSFGJIZIu3hUjTmzS2EVsfm
Rj8VO45H/Z9x77VrfJ8427uWV5SrF+dbCBRi1QoQsdVXk/U8dokpX55JifHHoTYK
f1UxzDlwTogdcP4uwdKUuPpM5y9aRsS+aCQf0xcW7r0jTTdnOzqAnL5LN/pdPM0p
BCHhfyZ6ShyynlHkYtZGg4H008/O5xoj5P2Dm4YxGL3zyHP8hHK7Gvu54+6oKJ2X
mD/LmrjKcZFS3oZW35cEg7g46953LcwScvReZbW6JbEchCD2qoAZ2yhSSg1QelED
NDCvKM9jlkMpyTtQCNzMdMW+KGef3aaDauFK/d/fLWljEddJ0TDW5bbCUbhJhmWJ
w2HobDpvchXewIXuD+BKLXf39Ci5v1vtz77pH/PV3wBtQUOczTl7LEnHmLqpDgrg
7UFmekCdLoWTHq2b6ipae7j37DdhdJ95R8mdqvoKREGDti+fuSOury1P2SPqjaY0
SNuz+4iTC8AKdCAt/xctsxR32O/KdHTGXex5DFOUf3fspZm7ftfvit6SpNCnxNan
O73YPqSWpFuFjbTp+jsZIYRZVYtqURNJyeCFjbu2QQfKbepUu6hooYB0t1oPRZve
qVmPmmjsyG8POyOcLykvc0bwoBmqto3i3SNrGe1/Wg0Kyj8A4I5QGcpVApI1YKT8
AkVH4O2G94/4IdZDfzNVko1+nBDJWNEZmRAKZ2BAlsCTg7JfICK+1DNQE8+2oKKB
0JwfZJC/iDLBY+nEwpcyGmuHRYaVGYUVlj5VF8FBSoFhwoNV38Ur7NnNdRgbnFqO
KiLHShUDn3DdwLxAen/B5nv7oxAMWGWI8q7ABeCbAOz3osJ0tGskyiJRVRMwihVo
aXTXjxbS7QQlUInLKLOE1/WGo7XaH4Yi6P/NTBQ6F2EIB4pWIjqi9EeRBddNnFzu
+Y5U8bMloiyAexZlNAi9Hx59+LpNJtgQX2CFn/c2rOePL6daOHmOplJn3SA8CZ0S
vaJKmBcvLRax6P/9AaC/IP2XpeDchk0qSib9/vkIgIJj/Q/qb9Rk4rSqTKTGlJpq
HI7vnczz6slxPqecVoOjAIjHXaLHKbaf/hs91wR4Ba1mUt/dp9UNZ88hWBHzTTk2
08+7q0ohcMOXpIWjUSPN+MPhqGWtrlYnjFmwE88GYIqpzwCR9eoQ9y5uhHCHb4c0
vR4GpEZyWyGZofibF5FX9u52cSSHwAlm3vf0+x4MwEMsCXiHs4jlfiY0LCe24B9O
dtFikMfSA5x3rAa69n2OmHI9Vj3mHomUf/b6HgScCs2mzqJ7PXSD2qhcEIesUprE
g2v7xI/pRkmam7EYJPOpbthfDDJcFEVTzN+Dm7ZmubEljadixUk+eYQ1KWtqY4pe
/lQM1x9c6eeu2vI0WvKEfH/k0r7wlk53X/M0/8WbaIQrFzdXucEdaZNmuunfbyEq
/MdU1s0dxFdpgLz0pZGg3gDGOCRiR1w1y2bC4CooPkOgh4zsBD3LPeWOSEos1R6i
YwSfj7djY3aRJDRXE3lXqDAhz+ZQ9CSChCG/WUatU+yzB8nZ1Vf32+lg1C7tbz0o
lWKVmomCm81bDsu6nvCvxufWtWFrXSI0vC1AmdW1AmWsxmp7/hNLwzQ18Kth147B
DtXSuB5+MN9hmpox0OPwUmFPuwHqDsn+Sy2tmE+oOCXx/vZ+7AtF9rtrbsNG1+Gy
0oOo+49W2VKm7KaYegDTku37ooWIS5/Sheqr+MppBloKvcCONN0i2L+xRZmDLg1y
1PS7pIP/vYtJFAV41ZCv/VcqwAGBIxLDeavb9WjO//ULCONhNFtpK5ZGv1rORnM1
p8R/ed8Wmp7UerAU8XeyALDUkkVdTWhgDTt5y9gS9zCxiNfsbgXIk6eoZfuTkPNP
9grLhpCzenzHc3HPkMTUXl8fAGp7IsPzAZYiDXjFGT7MtbM9KAT98fgOrHtvXJvP
Xg6HJuEruzFO/GRvRis1FOp0mKlqLtdU6D2bfzoytXChpYLeI66nXxFA8OAd5WX5
EUJauyNhPVoqQKjLKkuCa49BruW7b5/wblJR7EFo5bPe2FeuC9ApQrNb57yMQaOe
INIga3qWjpEgxKyiXliveJT73lpisqcaHmP2SYV874bNGAA1OsWocx8sJjjeGizi
31MQ4BflcgMfyLHKqpm+GOMFkJkyLHTGiHpt/kxDxCViHdyaF137EWvvKWQZ7a2S
V28gNGv2CctzoA7nzEnv0IVgsTRXPkc540Q842GvFPefFsckm+i7X2LYuNCQW6qE
akzA7/3cIOlitJSXOYXUWn7BFjD4BYJ8EzGzKvESffdxITr8t7dhDtgjfDxITf6o
HK89tY4dQsSmStrLxnPP1IQ3gOP77046HEjnKSlHNtylcjaezY6zUOCoxs9h3nks
xWElG2buk62nHBsVfKlm1DpuDS4N2f7DMjZUClJW+fzz19+MUzdRjsGk71QQ6/mL
XGk5WXU9NIgRZcQIqL5EcWjfTTzhsYxUr1SPzDYCGrlNt+h15zHZZ6tmrye7kKN7
/t5JqYRzi9mzFSl0q10XHZ+KDvK66rnZh6iO5EnxtEMwa0nZKYxpNpNnGZ4dEYO/
DyQImPIyoXme/s/gxvcg7wmCCO7uTjxDY8ZqNmB0L2t+4NyTQzgwZVz5uE2l2Ift
NdjKSX+wG86TuKyFj4Gs8p7Qx5oaMLKZRtMDpgWr/YTefvnzkDyGefk4JJihq1zR
JWdGY6QQhlADI+fSqZvP2UflA0cWCX7t4/dwU/b6mIcRyydVk1feThT4D1CXcLaA
BZ0WwZlHrlfwdAzj+snYMgy2ZsaXhA3D2PgQ0ZHqv0ZsxDrF7NVdm7cgKMlCnFAj
3oTBSD4OkAoA5KefiRXHYwH9OzEOmzADc+9o5g4aqygc6pgMOCzL4ZLJbIHtk4e+
0ajezumuG18Nb0Mr7sqxmtgAduAYI7YsTupl/6CVpIpvnGOPwuC4LY3NaXLRdvtO
f8S+wPEjDt9IzQcrziEgyRHBCW92TXdoPOBU563qp2cM325Wdt99HOZZxkrgbMoZ
QgUzrOBERZJhQTepM6fA8Lo7ZY5tzxzws8GvHUPiCr4kW30LzkdiBJzPp/NgErZW
KR1FMOAjpVOmF+rhR/KE9pEZXO91Kfv3cV3tBRzNcaICcznXh+Hlpp98WpGX5yKR
tyF/2Mo53lAYJQNXfYHpdCvhibvp9dcgWl3I7gU2vpDfY8U/+qD19ElQYgHpZ6+1
kzz8nQZfLgKY+Idqz1YMJDqiyA6iOjVLODCTVgEKaR5d0W844oLCgLbc1UbTv+wE
A9ZM9oktoy3RPkGAMM6SkMcRZDHbn1McVCUMmLQVDl63hdkWWwu+YxbX29KqLWq5
vTAU0M7wloL7nqg8OWkcQggM4Af26SZZ1J13R6wcuY/hJL0cUdY5MfdbU3d0NwGr
xw3z/N7gqqR5gqPBnM4HILHuwspuEK7lM10FUxIMtvMWSLnrStWI8w5hi8lF2LOp
v0p5ZOaAQB3usTs2FS6Xx/n96FdknjhwS8hmjLUjvYooIZ0HOxfj+vuPcDY+3ke/
zDK4EJIBofEYiM4HloyRaE+a2yevIvAXgEZfafQ492wfqnk4GkkGtqa2lkusigKN
4GBCC1IDMWda/j52DtOOUOijIrpoFwVDik5X+hBC8eG0tWkeQFoXdr3lRgGq7Qfd
jw8Dhn4XusQ1vDjity0kVl2geafkicsK4zbqOkX8b/9gWKmBAMiQBdP2fSAu+JiZ
l2XBjqIEQc+PFrp+Qbd3/DiCFbY/1aiUpof5+NBMmb05lUapzBJLsrzcP1gyoWtp
EXz9cj+vXN8l/1oMSHrG+9B+YrmmOAkc0x8k6mHKjrNbQkXVc5a2lCeW9zcHk1qu
S7RNXCTtKtFmCbwBwyFMnGilAICtDskwYv4hzqzASLb7/lhZR9FrWWI/TPG/rdvu
FRDQGTYoMDWuuPugB8rTRZUQGdCZ1eZm1/7CRmr/ANGd4KH2YglkchxdWaWQeJ2F
ejIJo06Y9wOv/oj2zMszPq0FLsRVNQBO5QvjH9o1tG8YOCICOqlJoxU895Kq0sxj
GGcnp87ZE9pn1Da/eLqSoA+bH5fjRAw+gq9ljvNJOCEoVybp0++H54yFUj0P+29Q
iJxjXC6qW++7Er0ekpaAy80evbhokdWwBkYFSTzNxQnKvKCt09oggYsxhy8eoFTN
ShhrsQW88rUq7IgCn+hW7gNMCOtIk9Y2iX+6lDvT7Wmr/lWf5xSw5NzFxiWzJ8MM
zCi5hzRRUFdrrqDIWdQn+0ys/4ItwY6gmj+vk87evEW4bsRaN260qnnBifGxTym4
hZHlp5kWYoptl+1J/x+/1z1Z4/Z4MZC0yAyRamijNG3UZiCBi/InUrZ8aQxwJxOl
2aLn8w/Ewz9coZJt6BhkiUJ/Bpa1pC/Uh64VfEZzDqzvYc87iGpwyildCRjT6APe
rxNFuiVtepR7WpV2DEzUbRqMyiBal6fSytndxxzTc/J1k1wQ5YulWg8O3sV4vGf3
Bu42IcYhrFQ9NRxp4Ripld8l8D2IpW8JS/2l1zE5LT6XA081r/Nz4Fu6PbSmtoBN
oU8kEdKMWvpLJZKu/w7Efk9RooM565LMS5p7pIgSt18zar8mB3zoWwzDR5esGVvk
fUCC7HgIVlmOgnwJvff+KgKhIG0l/Pg3xRvn4YLvPU8UVAsI7sRhBG8/dmackVnF
l8s+BvzonZk3FTUETeICUETDEoiEFyYBGlwCI0vwCR1VbOH8B4RC7UZfvYDwXeig
XbSiGaf1of2DYPHl2ym0F3J3o3MdnjJ+Yek7ZqVHf/aNzEXn1xz81cvx6loC5Exz
t/OvyZD2hhcUXGXF43UVSSTKRmai8FpG7vafg91A7QzVMDs8Bgm2Xe37t4joMWIk
ufCyxBnhe2p4VO5aYt6a10vvKR1ftZQEpP4trTOPGf+o183QK0e/JERCXSIqN5Yt
UadDiaOCgblA/iXQ+r4myTsqYNdPil3dIgMe/62eloOhykyoOiaCgtvkk7cDG6kt
By/cD7P5Tzph/qtUZOFqE1mIHY+tYPYYKCxIcS4pLiXfNaeXGFXd+phFWlIvy8lE
G4u/r+oRwIkYHLz/47kKu32L7rffxUDBkiCdJbygPomeNz2+M/9tX/vTEfDiNev4
XEMyK1+Hjp//HENmHItk/0Sf8YbLGib2m1ae25Uu8qyYztd+tdKQnmU0GPgj4K5R
wp0aQ/AFExAqoDIK0rluj297fwg5aUEUo5bJKDwZXKaRuvMnNoWD5jW9AbTWhBsP
xQIsTIOY/PIGOzaqusQM9xgknWgGodgZ1mlnAzzIu35r26mdjGbejrmGd67n1QsG
EU1QbBYW0zS2tNWA6LQde3kH9bS3umvFAN2GN02b4Fjvl6RoNfsNMNmnvwPjJI9B
uOHhlVtGrrwVUOjAsy2jX5OCyHFOjXY70pXirSIp4WewpUS0YKixh8aKLc+Mbxm0
8sqmI5+CUKjv5Snra/vk4mPFKFRHjFVcsu98zdJQAZTZpeGXZe8bKV6KjU3l/YGH
GDO2qCTfP2JvVO0RAJ9ofd9Sg+Wmd//ypH5ipDQVa+W9pQw7QCp7M4b3A8jSEklb
sxWJdryiYZ07k7gfCyClRlOcB2vOv5Khmrdx17j6akVwjiCPLoC2Oqz4iuoFmDRZ
TE1NlU+PBqe8cqAQonJW5SCsXjxnN/tcejJhrIcd/mVjjfG5WA2Rft/z+usbVwM+
sxRIcxfdDtPHtgRXG9nJaRKWxRnLPQfq7wlIlQw6DAO/+2yYq8OWYjL7BRp8b3sl
ioYEAdtA4hX2nJ/7ZhVaJL71k1o7C0E05R0+yF2iLBvW79FHb9Nge3KfvSE/Z4b/
t/95WKs8lHDjHDzSNGFxBC0wGrI3R9WD9b9/j0fRi3gPSZoBaJAtXrB+4uFDG8kF
KNpFAEnkJgQI87gcCE4SetwdKwxaHcyrRG0olCdgmO5yz2gHGQ+1mjJHYS8DmvKm
wai7oq0s5+yDISKMwxtRVl7d92tmh1zeiDacjCZu32qUUHbIlhswJ7eCpsfD+v69
I2W/v3lEX/EpqQNpHtkjPgkPoqfYAdeVVz++4cSNIgPLr88zltq0SUZaQgC+86Y9
Tu8A5xcxN12u/lcRQnKf+N/h81iCkQQ5ZNZZ5dKI7VzHU/6Mi6AKkt+wLACnwgRp
cKZyZ8PCvD2xhQ/Cm1KN64xu8UWbe85F6gW1DFOsuqh/jkHgCWTUe2YlPwbckzj6
Y7d80BEqtKfUsRJmmXXN34+DVKzJw2pNIUq1bPd5GWgDdnSVocLxjMUe5gWasTNq
YTtwHMBSAPYpBItcRbzQ/cCOER2Oh+w8L6AiAq7kTjhKLu+cogq00eIDOn7WS+B+
LHMHiekSxWKYeXLRVlgIUJ5Xym5piBPWYKkfMGbMe/BVzj32Bq/EGvDEDIAveC7e
RZda4E4gYh11xX6nBBYf816bwPUhqFG3kt+8Q9eIgSZUcfs/ntRQwGegFF05lAOY
FrKNND/kwkIC86HaqNlfsnohImozK4ptBjy2r0NAAXBJSmjFPSiMMoBs2Cbnpey1
olzGKVJ89YVp4QQbbkNwTjAoPxSxvol3V68kSgjzFXDb4CaUftURvI5spniifTWK
ZbbmDR+ikifzcSXn/K95VtzoIz9kyRd5OySqNc4RI3aeAk5qoVEW84yTxT0tNzJn
RFv8fZdK5kX5tb7tr0U9BEegNpiZuG2Bj7F9Mc3aZ8NCv34AyOQ3NNNdjlgl4fev
PzKssyBnQzKHuvozxx78tRIEGLrtUeYucnQAjMpPXXFdS+lLaEUTuhHxFZvCE55G
tVDRWRNnJiOWP/KV6SvwPpD0FLqDIT3Wob9HbQOZSyZTlEAIrbNfGOSZ1rUyV58g
LVGwoAkBhhYgfmUdT/IlHqaZKejxbMpazLw+SsgzVxHCrNeDdWncYHK5cThsidif
/IPT8PqdeyLocIHoYpvperL2xKdB1m7DTmH5AAEzDgGcAzR+tjjlIlgkH/8ckJnL
752sQzP0OJgSw/7tH8PO6dAdXaPx1zzN7cf8wCJwqYfrMk3iOn5rMa/OV8nNVzgM
F/R/Tnbg4OiMIvQGG5LVm2NgNiNvsI42I1n+DXaLfomWYe1uw4JVeFWRVxhurBd5
SV6Gu0ihh3MyNU8afEs3KPq6xvvsSPnN8AaU4ivGtku7Ovg2qgSQ3u5U8+HslqM0
Fc6ovsgpFXiTxeb8c8LRQ0mLl37PNQPx+sv37WomWQqathPdLzQSy09IaHPE7bqz
yVNWaTEwxa+zt+3k+Cn2e6VugwsPzlnEBlpyLZIY6YwDozlDbl3ARzq8OmILVldG
c7Y9waYWYzQ8b9QqcD8n9sQqldV9thz/+zQTemO7W2qWU7AI43sJHX9gP8e/WRF0
vmhPwht98ZZupgfkx4liKIxcXzMVoG5UItO5PZAZaSoLHpkFLxj7Tx57NkQ4Dmil
GfVEV5G1p5Ao5RACqI54FOxMhL4fwqT89YibSaxSwOEB2b/DDtdi5x9Vqi8kCvU4
/V5lCIf3k+6lZY4I2Qz3SjUoPKa1mosHyOPGOJVy2S4Q1yZpmW+IDJ0Nv8WSMBQ0
A+IshtQ5+41dNWgHN9QPcKaRHsLQiQuMRLVv+gt06PMWw9Sh1h0UXPTkGFvvL0O2
UFN15Dcr7Lt5mB2FmzBv2JrUbTJ6mA9oM1inii6gJKDLZ1OP40VlnXof3VNUw1S1
wfAyM+q1P4nOPGnNZJZUf6lI7UlbqxLPYWbmt4TmvsLbvibz/VIP36NWB1mmrjnV
3+fz1LuaAlndX2iQZ4WmDBs3kZqAHaZKXQxt3JG+bItQwWN+I3aUDtKHcYMXFVP0
gMI6/v5CapcGW9DZH0Qz/6Q3Pj8sKdAy5cw0nAAHX+P3yPn8E0TJGlFGwoQ4g3rp
ev3egrR2wOImXbQKkEd1hlLy/Vb7Ki/+iS7qJaJEmJxoDYDh6qbMrg054Ji/eiY1
UefZJH6JEUpUf369MWY/kohehWfHYVgn0k/jsekvrFMGYa5RPZ955jm4ML6cvG1i
wIPyyBctgQ0rpp6ZrapVIFaMrve5HZSSOfh+3CuP/x49xXOH7yCP2O/0D6LBmGxg
2+7V+LygZ15lGJWlYy2xOp2/eUgXWG/p7LNAvWJPU526aZCfyJs3NmsHKAJfYbJV
SiKvmFIq5MO2iZPlqmLQ2+nexflhcWFs3f90su0+qmLioCuPaWa7P4JGS6+ItHiv
1TyAXH6Rm5QEyK5y3/tGR+c5vR0X/IqBTNuex72B8p00z74u0zh9dvtAgy2K6YaK
Kf+RrjoGoorppyAVL+RqghhVQTxXdiUSmQvqnsTahUK4cWnmJhlmxnHRGPCxKed2
TTgTGcvG0uYU4QgUe2TV/rEogQThU2FiqdY45iNOejswZZL1vL0oBgTRjbiSA3++
gBpIiWgxGCT8d3Uno5rLIdEYVmGf+xj39TThqbLuvU0FAoeyXwHwoDyseA6a1TiH
oz4ewV08QbUgxHSdZr3EY+MZi9iPDPcsd08H9YSmt0UQplxvL+GPNBJopuMmcO5W
C3ZS30o4jPg1wiRkrtz2XYZrReUG6wRdVbFDpyUXsWTYdlih+bbcXGT8jQk+staF
TA9EWQu5EPMTrs+Ipb+lO9hG26iJSTRtXyGsYeZiH2vehXEewRvB+I9YX/eIa08l
mzgw1JjbQkppT1a59VKNHmlS8OlAA+jV0GAnAPDscnVSk1Gn/X0iqkuyhgq8/sBb
gy7YR+RcTeg3/f8iUKFIwYTZJ04F4Q02ig4Ku1MqA3jn/eT30FywvGG5cErU3xUV
5Ng/sD6UGOkZjCV/5Xvmgl6ExwPcWZw8e95T1NyD2+Rsg3Ra5B4MU9lu9Drb0uO5
YIMnkrAj2lwPWYkRDCo3DqTMBiERPMtQkqtp/rLxbgkxnV4sRjpM+fpCEdMbrD/q
mtLoPyxWsIlqrA93k77l2K0KIkZ6XJoqTXedBnULqVHbETZgZOS+C6TmHF2L2HoW
wG54SVgl3HzPX+TMnqmMmGmefQCtUI23vyN4QBe5eElkCBqCRs60CfY1w5N6k3+B
2v9m0Ckl7SUOtFdLqiyLLOQIchsUp8VWjazqvE7dYc4viOxRXRCSrOKepxJyZw08
6ICwWVsBSCE9YAjOs+6L3uTRYjsV3KZqu02ehMhtIffXZm9nOWuN2MF0xGBZcuQh
PaQAcJVkQZqE7yqhBMwdhFPJDckcwoCikRq1SKuCVTu4g2JYRiJ+sd1xvLxX6e5c
LWtZf1IifSUDtr6Gg4jiilP19mZf8CfkPvnmt9paNtsM9Ltahr62CZgsGKLAmBOb
v9un61JrK7RbmuJp9aVjMpEipuremzT/ULWpzknJKv/srk/J87gsFAQgpYRmJrKo
1zBVNVWWDXUp4ThkhaHNv+1RQ1oaE2Wsa8N9g1OS9nao6tWNyYd5/EvVANKTrPnp
GAufLLzWLSmnUPNkLyw7qSjL//P/OZSrur/ykkLW/bh0pe9fGn4E+HFlQPHI6kLD
jTO92heIO7GOH9ZuCsHh/19Oer70nosHEnSmvbowy/8/7Azxr0C/paRjTk795sZD
3zt/wK6rkzh86HB1sp63Z+YIn92SPDl/8jrNBXL93vVMkDymKWXNK6He5zOq+WBa
dcw0cHWApN5YRLLsNmQXJvefW632avv+Y0b37PzNV45CyPLYs07VSrm3gDvRpyXi
daZUlVVZlyNoCLuS9iyAFg82DS+8+m2oOnY02IHm0Q2w6br8sULINyhrEiTfMMnU
IWAb5kIoM6WFchGrGAuE2p0nwcq+UVC2PrTXJrZG+P8uAodV7f5tFqZKFVW95Ib0
pwsGdbKJhCCwYwWfYx6so+AjW7N/M7rUFqC/0Qr5kgDJBgcW5GmscSBXq0M3VZPq
iOe2QofPqxw4TG73H0zeiTwxAST4jCZBqPgdBvqlyaVuA96Hjx8pxqmmJvY8mgIb
Oj5eoXuDPnjMTo+RYjoIK677hqtbsdWfWbvIhPnCtjOnvH9Gm9gStvDwKBstfpTZ
PDxK/BBQxBFCmDBZo3+FJbW4Fre7+0xtHDO2pf8srt/sDPkL1no2n3tlucqdupLz
D0dsmWcCKv+2h2/Oj0i7uly/jKkS4axCvXkXF79mWc0zEXzauS6PWPgzMsuRC2cI
WcQe/oLFUgFu1JYIozvHk7JtKH2HaBhNLmx6w9iNXs/CVE4CpWLAAXf/xGQWRsKv
Or5bXQ1rJWTQB1fOeUuD11P4KiVEC0iF+tzUl5pW0LlyW1t1ajN/hogJWvW5Fha7
Vh/QijWIMdKFyCUP49jNFdaHvVognA3OixDbgIHAmyIxUA0bM+d5qdOIUp3vBMbk
PBcZk8t6hyV9+AA1WSKUVGmU8LFio333QiIpZcVUDz4bDwlriDX5qpfpr/cZXe5/
2uIIs9jJHtlWOfQyIGBc692reyzWUKBizMsmS8vf75hB41JBR0ECiyYhdzrcMHPT
vR8T4zqFddx92mUJcm0RDfW8PfphOoW2MiO/avdHEBmnMecedl8PRoIkXgbO4bG/
5MU0bYVktljk9p1HlDwGEB28LWdmXh3oW9BzutTULITc1ry65F62az42KfKo0lgE
KnxZCdsraEjUeHVDd5QkUCruITzMEbaLuWqTlZCsxz0BvY92Dt2lX81UtvXaqtN6
9bHjxaqckBKEWcALXl17FiDf+WbApuG5gXQrnra/CWF0HweHjGZ2ZZNS1w8z9N3C
WvgrA1/vu131DoqYnPDJtfgK/Fqwqv0iQ+k4kXATT7TzGREZNYSQrxAVJndsmgsL
9kjwbmdA9dVZQSdHPYBwfGvrzb+9pZfltDw7lMBmPn+AlZRVc0cv6O76D/Px+wX4
IjT2tJLT7EX8R+pFU8nELS+fJCXKBwYgCW5QONF1hbtQ/xf5dG4z8XGD2IOLGHPB
65LVtLVMi6RwT9lt2eaAGkF09UraYlEved8ryCOoTboEMEwQp159iyE+Tje1h0El
icXsQw+ujJF65KVajfHdlTPDQglAqOCtS3tPVyP0P9BbeTWFfMDJHThT6RIKUBHH
KZnjHg6V36o8tIvEEMpP6VsVPp4sf0oQ1BuI2vIOkpYX+dGxy/G82AqDhwWh4eWt
oiDxaOQx0sCpZmu9jMwcGR8TzexcGSNeMxA+hJOQdQrbHEW5wPfE6yNh6b1chQ00
yrccRIG6oI756eprG08jg5YGDpl+vMNI5S6xPgeWRcmhh/Bye7Ih5fQAwLl/jwAX
3/tbz2mucRnF23gZt/g/xgvwmcNc1pQDcHjDnhLGML9aSrILChUDKl5mEiHdVkX1
cffMLT20K4Fcgj2Ai7A62tU/WXZTjm+SrKWa0snHbE1hKVkKXh73AiGy5/oPVlmj
TNqtW9o+TgzO7gihlgVMTuteWIyk9u1Pihrwm1u1DqLI0yfkbyqoAofS/pS8pyk3
YsDqwt3nxcTxKazWhxWvrDN4OEc/wIb7MJHgoEj2pgA1MBlVmp58ctqQqCks1QAr
FApnFPoZ5PNBL4CqCNxcSMivTnUVBOAYZV9buVFjWScQ8qFHmy+rNefCnH2uvBlj
mOkfFWAwvcaT5IGPUZEBT06EWKpE7CV1LyIQuVq0xKKJDALaiEHVKoHGZ/BQdNmf
QYPRYC/b32Oq9D/V+jPEj7GfrJisdhuamCrq+8H9PEVrh7n7YhBFpiqtJIIzWtxQ
5VVDMQLGKgbJlawqQXuTg+arOiFSYjxgBQW9ekK2aZzwZuccCBTRU/sRTi/OOiRZ
Dntmpatyr+d7qOod7DWPiHaQfOvfcptTkJjoOrSKBAS8XHsRfMc+0d0GjRWs4w6y
y5j7vf80Ljh0v3Cec/PIgj4/fVCcMfj/ERPpNHd72tF1EHr5X8z2cjuE6mREF95i
Gd9XSarHf4b/vICN84BtGJbkM77HAuAASVkCWvdRKOpfBWPox9bJpu+VbSu+xEdJ
Qlk3P/CqPzysm4FV2ChvD53ZWo322Tx2HaM4/DbHq/dyKELyJJBLMdepIaayhEL4
8cFK2NA/Qbcl5+DVhG3hTQZFtxaDW3RvJFToeF9WQnMjJkQ2wDCIaZra1wr8wBCM
jOGfvmCDcQgaCs/2Lo/SWoX5xbpmlYRQRpINEJvyz7a4Vs7nh9tU+/uwXqUN6I98
msNEd5vzK6rAD4ByNhF59wdOVRi7nrNBHB/PevZJotIhQRb3MvHmvYSm6LMXiw09
N6S/57XBw8S+85+o4Fvn/e6i5RXP9xGp6tbDACrYgtIDQbWLlHZCh49N13ayhZRF
7pL607W/5KaED3LirdHbpZQQQXXmecl9k3WCff1Y19fRJx0GNlTcAiaCvJnyv36n
X3MhKGDEE7YJm3D2Yz3CMKvm+mFRTci8saippEWRLqnhJ9UZTvTGuNv27W4VcZW3
LQkcjQAM/BZ4K4kUTSUzLyNO8Qz9o5uj0Kj1PbGKWAQmrNq55GcUuh0lJjoGhp9s
0ye7rMXVv1PH7bAvsEvB6pFVpktm+NIIGVpXR1Z4rhVTghAopz9aAr8cPlDgFzN5
nSANRIuf+Srzx4VmQ/hzV+OmoagcstCjOTIsvR/abXbw58rCsicoog+qWGFTOvxs
+OJMh0x4BGwy4yMdOTkzuZaXVu/zslu/5YbB3lRfaswfaEEPMTfgUMuQBVQOI93u
dGyCrGaPc+MlNLidJzK1mxPr/yRsCxR6kbm887YzDKvF/5rJU2x84HNyIQh4knGb
jV8B895+Zear+B7aa8pV8r4bYOtUHJXMhu/kMUKoyRwZ34Oe+X+ncAkGznOcx5vf
t3J4obqqCdjUq3oivAMMADXtkncsbh7Ycw2BTg7ScnyqBL/l4kV9IxDRZ0zAgwO+
egob7y3r4b3aqpqqaz5G5+LXIXxtPTwnAFSHb32w/K9roRJqGCX+V3j6IOUttVZ0
XfHRmav/ruHidmdTuw+5WPuBF0kzYgeqCBl9kDMaNNANVZ2NoKAAKni8/ZpYxdSE
kRjyn2N9KDGtgxlwHVEeUBhTX+RufxSklOl170G4RkKmHs7ryeztBui54cqzwrDm
D6KSN33N6xzeEAs0EbxEQGWBz78RiuXjDiORXUMTBuCYeaQLmyNF0/+rGkC2DlwA
OtQdqGwljAKunPHNORuhGbE6wyVgUgbd4zn6iiPNTgRu16ZGBWkhXbprl9C4qVFI
7eArjmdWjDa95lA7qjsCw45NYZLhGMQtJnSUd8oVq7rih8kAd91a6hOHuV1slgE3
Ql9ds5zavLXX8E5AvG7IE5IIaf9CSeBLqLMVukygX0s9IkoVsqH7KoddD3k6b2wa
T4VbvPYyGluKzs52nYxqySCVYXmMkiYkAoa/toHS1JuXA3GNUczsu8sHIzuttRHZ
7kupuwbx/f4z3AZ8q1SES1RHpmzNZB2Ig/aAzB2nwsBBWdGBKphNDH4zQGv8Pxi5
TeTULXiU69F31ygtDWxTxt04yS+iSH3rtwnzbJNllETZ8LuzhVjK/P93r2u5rXU5
ss8D9Ds1Xt25kX5w4gLD00FXH+WqDR8uZZMrNW8rGvKQ7QSHVVXW1H11tajyMdI5
pCpGrJby95g1Z213qNXnQanuMDmyJ95MgkkAZcASEqHoCrpP3JJGmwkUzPonZfpB
44zxWZH2v0lbUA2VUgoBEI5hPDzF0XSJrV/BRGHQdKV0ddbWsDxWEqy5lA8qE/lX
txMnxJOGCwV0wbexCeMR0N8GO5u2zSTXBoUDxTse+TXeAfF6bNnUqAm+FnlZMlLm
92ycuGxtZcKoJu5SkRrHJW3h5Yuo3DMMc3R/8vDKEcgxX4cAlzxjwr9SMwe9BUzg
TqJozYamKPYEuGASYMTKOvujUDlLtX16OTf/KHvaMalpQZc7aIEgzvg/H98TBUSR
QlTWm2DleHi1SyleA/yO7CFXH3MQoDrErxP9cSnS11ch17NyM1ZFX/1SgdPJVQGU
NVA1AGMZp5/bvKAx4u3z60wAJRyxtApJpr0/gmwr1bx1X+fBWbHETlsAVmlmAcfu
maIkMfwDVrk5zH8aHvs48OinyAVg0XY7EbRiHRdhavpa03SIpU6vctKsLfdSAWmE
hue+MOVMyYT3WtC5tna8X1iXCMBdzMokiomEYZN8YYtyba1I2WavWoA/4nmnbPgn
ujdSP/eexOS0fTel8zmZXMVdKFqXo9rs7cxL2GAXO41BfdCqPMWXtHnd+Pwzq8jk
xzhSB/EB2myfEvMTC3lIUpFHqlIJeQBaAhvoNh6mJFTjXuMAPHqe2VAcQdSANzbf
0WuDiN4ctwbvRQqHDe6kWfmLmN9SPyN4MYsQ2F/lZM1onD+cxf84pg1BMMMTh8DC
vtsCtKKmhoUV6GgpCB4nXVMi7pEeZQxAooHt1rVIHqaru411jCXAK6A3qyt/EUT6
jsOZATOhc96RJv5G42R16O5cGF3CK8iwsuy9xG9vjarmG9LIQC17kg4o5Z3317lI
FcvakfkEKvm3q/bpQIyA4gxyBQWxBeTCegtv4JE5DwXDm09YfHDIO2BcpH5gBPQ9
RPqEMANz3f6M/CvIk9NdLDYEbhlCWXc74pLZq+mruqB6myEyKpsvEy5zpqhOf6+O
NQnxpXlugCLusAbOpXSxI894vTQgC2tqwHRAhpDhVapC3T4hqLFTJlU944XMfrpw
qfJsexK5JZnapZTkJlDK6TiLp4YUQ0r4fYUqSLGmr9qKk1G+Klu8zBnQsZ+IHKDN
QAUHMWu+Dv0+gAUjFAR+kp5/H8dG+gR30CwqztYD8CxPlq1C0hgznW5/QjgI+yC6
aNgWmPUQyuwqJEGChLgCZxVtjwSKaNRl2TmKP7X/dudbnOdAYzGXY3g9euySP/S+
yZ09JRbwQyEh6f66GmyjVSgrlc1HcrBvLn2G3dJ3FJS+SfuITj1brESuexX2RTDN
1DCom++I6Fmm9u3HsjsXcJ46PLdmwxRbXscWMP5+5ah4iiCOgIyy1sxlmGOQie+b
DrjFhLeFb9O8T9rfHik+AZTs//HKj6/b82uLbQ2W0JKmgbUcOsVCEWc58LnrQhcR
iU7vzvLxJ7YitUb5U+p4lNfPSIxNWHUQlv4iiw7M1shB6VSzAyz49p6ievkH255k
w8i9d4OJTiRAgjKFr2huOTIJOWvIRgFNxhJu5SnDRX6j7tjCUkx2LoyIX0haaI2K
dPDPuyzsEAcXNKZh2KMqIhthEeye33gfZLo2vgevN/Y1be2vJoI7FQIx9YvOw6rM
cUGn7zetyLXLXTvqOhQn+k8TfZqVQK/GvHwrHIAFMPOrqqRxXytbpCHpPish3gRc
aOe4sm/028z/Gtnp3mWF9CiBjEmL9aRKiAjN/5etMh9OKGkUanOVqkCgyzJIC/P/
rsvg0ykCOxljinPt0qCseoI+1TpXTfVaa4/Wn+EjukxSYkw+LAN1VnyP3AVRGy3m
Q7xaslbTB++GLpfmRvGmlCL/6oJRuLkPyWZAVVaAGUZCI+hoQ23pcmyM2S6w7IQn
dt71FPQ4qlkhK5H9jXwaYfSLmFwthGnYuuoTi4sEimL1dYeIHEGvrVkEbfMwYv/T
Z/5TXjX7yFy2ObogXJQaQteEZteD6oK9Gus3H/VZ2dXmNiymAKqSD1ZS+Rb9VdDu
WF4sRHZJ4Wj+nmoGPUWogFpRIO6hsqCD9PIsClGFrKk9KPy7Yn3pOptnEJxGDV20
m+J0Xi23jX7OhbXAM2gkWirZ5OZMLFT7OGUc6ZVy05tbGW7f5F79BpIMBCFqF6tC
TibxTGWM/Eniaj5aRdMUxeAYSouQViFaQXpweqvazrtzbnSMkpISjSOsonqV5MLd
9E7+Rlmzezhn5lm9FVj2fRC8roz2Y8BFUlWyHYBOT7Gkb191pCmOL9Mmtfme4/li
Wv9DoBO10BpwBPkhsZVZhHMQC7xjogTWxEspSOE9hYk/47/7EPJVa+fakhC3ANXr
pfhgGORBu6K2Rx8PBq39WFKwRBuszC9uuCUJI41tXBFZOWqFDUBQx80GLlgLuLMZ
FTn0DlSxdky9rk9f1//kMqah6O6iRrj3T+ODoKFZ4SXt2QlqDYddzt3GMARDFqcN
9NG8V6k24p5w/MgrHbOhIi16ZmmvVUc8M+1pi+vkrRVdM7Y6QTF4JaXd75Ll23Da
OJacL/QBBr+d5akj9SzXPu6N8m8jEEQFTf4F8RbyOZmTFCiz/DiESBH4fV+5aQ4R
IvSRmtNEyVqMrwuALYmCmmsyj7s9fAdgZQ4IdzTDbS2JwQV/+DQrtGQ5ZRTaJ5GW
FWWR8UnRV5H0Pbv7vmWKESdXp9uAb6Jt8hBQqlQh095CiehO3e58mhJekvMmQ1/d
pXURZA9/dVvFNTBAB1IdnbquSlciyuX1YiCBIn5Hz8Twl5ntlELDMDa2B/HyXcqU
7/Rt7eXIMEOb7NjCYXqOdB6OASIe5rKGGQAOve8F+AY/rkaHB9xxp/rgeS7S97dI
G6mgFBnz5lWYUz0F3/4aJZiHeaQEn9sYGAVi1ryr3e+tFwIQTcoU96TYbuC2d8KC
yCpB7maMYs/ME3T4qBgs5+Qa1dBRFqCS5C+dPT5H/+SlOVoMRSOSZQd4Dyea9al3
WFJhGXBeaQnmR0nJ/I8wrizqXb+T1YQMmBui00HrFuayZbD14urmpi0IAC/b5TUC
xyvR4N7AHOidlkpV25LNvmjPghYPXVawBnxtaB7sibk/6lLWxZQ/X/ElpgB/2F1m
HAAdmn1R2q5CqDJPtLQa+9RSQXqDPQCeCGRZNdnbd+sGLlEs/jLmxwFkiXcE1ZvY
2Z00LZCDSs4oqVdprlfVUFhp+opQlfCEUTYcpjHyJRXiiiB1wBS6B+fTtR+REWDj
S4vGHrPCRQ8qax3AAr+O0MeCRLDrzOIj89cxWN2sck4UfETfuGSBamSd/xk7LgvE
lp8vvXS5OID6+lzXGKfQyLlIufs8vw7AQLiws9+V9d2BoLeOh+mv3m6MeFLF/VfS
qzqtGti7fMUEVKCTPIsUkG4uVE+FwBOtF9vS0n2G0eaP1RbeO4MdP22MtzYffxMq
d7dQ2WyZPfTKEUjLFzTdqVvNmbF4B8kKCJ1wr6TK4BtHXZUgRlmSe2VLXHdL8JxM
ZiHbspAhOAcMhDrV4YXQpnixrevvZfkoIEw4OmhQfp2OiezfnEW/RUuAI1dRakv4
iu+vYuYtLvGN3VvBzrWKIObcjaj5mBJyr/XXRQGMfoVrYZZ90gNE7ZqMm1K3uQqc
4Zmyz9ql84i6O9kmHCSm5VMQzU+HtcvbuDCCOeV4xnxrnarDZCsd9BlLX9HXDr9R
Qtyb2dT+i7HHqiLeN+EGvd+jCYEYBW0IptBETRIVrDVJAJJs/yqVq2z8VTLNVvJ8
7ZwADz5Vh5QnRzAYriiFWuA+HXYWukJVEol7i8GXrmh5k+k7AtwQOcPZostwcGcb
WJRnhdGjHjNfRB4i4jtStsjO3mbD7PSbyWvqip8cpaqadiB2nK20AkjYDMypgdwa
wBxKhxVFKFKdTnKxMeGVfKkaiagKnWcETHJ+SCD02q8L+a+acL9GirqL5LFF0CY2
+ZMS44SVS4i9f/zeSKf6pfN+EEG5NigMc0A75ZlUXSmmgTMGn+N2U76rlocaWmYB
wJB2ru4XU9/rk9I+0ygCDLx5aTeJ/URoNDmb+jPjdeiT2WR8bMHQ1GYWDPDOqP74
veyS88IGsuH1ZD3Wm+yQ8pBhK/8UXZ8fIRfHZ2QV0beJRxdH0GIlDVZxAGR0uXHM
op6dPnZkSKeECPH4EQAAFtGzmgiYvkMuX+ravqypLJa8I+wWp6Yxl+ujr7fLQBMt
BOVAg1GAdW0N+wWjbL5DX3tV/BhkKNoMPfcr17SYD/Kqfo6Yc57636v3MuX0R27d
0Xs4jpiMpTa2ok8a7qaKZT5fZaQlnpMLwYo/7s3vQ5ZhPX4w1QsSyHRfB9h90LgR
vdaWXpE1v6/y+j3MskOlOby8Koxoqo6L/JHda+ylEmcGJiFemWf2HYFOaGSytCnI
cZH6CINR3B+Wq2rHUyfb22EDo9jY+PN1+uTtHvYMMyslSE1qWeFmJO8V35xxw0IG
6RXj730iChQBjDn2hqEgy20FjiNXYsNSb5DMTpBFLhyJGJvggFEsD7W3XvoeRxtb
JTAASfZyypCX/hPhZZ+EwQhyoLWSYEd1OKTPjMQjz5UBW9UrERX2N/ADmPzk+7kO
2lQKFya5Aw5xkDWYEUI4OHjK8zQu49ZAp8N5hHw35Pa0OpnkB7IvOCUHLZxs6+8A
53MqKL1ieKu5lzrIDUrpQBVwn4HoB5nX58ulJy7wQlywMEOCWOAxGDi72TW0Ontg
Qd9R4KsZCf4JUFM52aQg7xWDdiWn7HtAh9/nQSKWbiceAqutV7U9I1OJaJorlWWr
gdjF5BbI3FyAiCzrmtYUDhyt5PfMURqYwM9VI7O2FrizQ/hUc9JSRmxQXQ/L2+PS
TZTXuZUhhFpW+urYRurzI0uX3Y0JEmHfT67M6XpVbfeial883dVgn4ITgq6nSms5
VRrr9HqE08RpG1KbtyXwRbPQwa2UsNo/zQlRTg30W2p9RwLRHEVkr2C5LEAjUNua
pvr1WiZq6d4dC+564g94V34VNGMhBC8ck+hfhHOyGvIIcL2D7nifc9a7zEvdVuuY
Ap2A3Xwf/Z94ZR26z8jisWh0PqDOAMCkrvX+cp82qwXVdl4E83VXaTXxZxA7qcFV
SSqdI75IZMDiCvmF3/Fakd2wyn2HOgIidcJ/3iMJHOYBKfqQUYg08ulCWpr11cVX
xwssZyiPgJZHqgnALUfmW9dB9ljBN4at1sydpB7KWjB3B94sfWY3SydBwVm3PjKC
xYA7tgK9LYS7iDoFMc9HgA1AJBqNavsDQBmQUXdohMQDMiMkR5zYmLXy3xlE/H6r
jwhxmgesgyGnn1ZrODU8VYez3eGPdxUtcWpM2C2+5Muf0ABR3cR/9HaUrmhfi73u
JzlwesZ6mj+6iqWeo5pNJdzTOQnpj1eqRQgPb2VmZ05k8+v67WVSebCsidLv4eqq
Eq5nMhLz8Nei2v6ljsb2K35M7+wY0Rrtnb8aMrVWDYJ3Y0VWK+rU+AmOIcrFv4bf
g6Oy/OrajHp2bNlk43r5E37AJMDGq50Q+c72mzZq87bugFe/2L1FQYGedgHjdhIG
Qf/+ix1DEgbvbGvqifQ3tAwoOn2xYLbGgfBmFiRKyo1By0afIgMzWiD36PnhOB/z
E2wYNDWeluET6MwISiC6sJ7bBNdVcfqjtMn/IGDKaf0vWgQyxfo/wGdx9adCytR4
t7t7AFo2jwY0Ev0Or0a5KlLueQUGpRlUlr0OKOXLrCmzSNKu2HYmDnsQu3nrwFrk
CFSKBE++3n4g7GOVUpM0tbmvWH7j1QJZW/YKihU/GUk37F1s76K7nbaO77K8lFVb
08Kj63TQYlvTkfo7ItbVQLYUGJJy39QhEmb0LRk3VCEZDGBW+EgkO8qi1f7MaJcu
0qYZ6cDXN0u66UTu5wqMln1/3JEv6gAWhr6GdK9m+Y0pvKafL/aF1UwKXdEv8Z2E
hlhTPT6R7+ZSeUK4BU3RPfXI5aaoSmN5Yn1lGtgOO0Ni/8qgm0nhSs/YgcG20QoA
SWwvCKZkkRqxmADs5zKl299hYkIkcrGtXvJopC2qcmLlZtj209WqjZRXdSp4yoiW
x8MDdS1E7M7zyBu8mQnlnpYYkfOmhMYMp6NJxFOxpORLYLtpac1QZOs/BIHiOcrL
7w6ZGpq4uvKEmqLScOkXKrmfNJjZmBRE+3/9QtNGU40H+r5ssH4C4YOKmSgUa1oN
u7CDw1gRAwgnJTBhPFCxib+BgIu9a0/dlRitI7leAyjDEwmlcZXI9AZ/GAAfPGqm
zaebyCvFVEfd0h9BhlGSHWCTpwitpr2Rbu8j/KEKYFjSrI1+vMWgYe5W2mUGvXIi
tnUrO4sjoDim2aZYMBjEocf0exz7cvsh3zdSOenKouJKvdbwK0pGbv4I+zFHbqa3
szv0mhS6h0aRrTJLiawr53fMsHulyOZAfweDA+3UoAOYTusNzJvDiBvb0e0YShUu
Fua9fMQJYapnaFVml8XwmW7xWnYxcbX0MpuYb1AM02QE/2U6wDnqvvuauZM+vPu3
Mb9RgjprqB2z7x6ZaAlRltx6OhPD10bB0rpaayfl5IlYIDskCD61tvINa+n0Rkuf
e3p2jyDo3hkyr+RPCqPUqzJDt9ysnfVRPyZbFmbi0FzOnFEosofFzW619DQ+3vJp
5eHN+7gjS9xQ4uhPZx0xsd4AMjwwUVoH2Fys+RfsLzJLLRBDv2u/OVnqjZFue62E
pnnYfhBZWK72vEPhmQb3TmXgOOML5fkWsILL81AGVXr9ge57zDdJvgRGxvanBBs1
BDGKZG8ERsIj5kTxXvfVTR1CYlkoe056+fn5hyl4rt+XRawdMcPqb7XxDdk+eW7C
9Ps9o7LiXIW/Gb4ODIlXIBT2H66SQzgca8Fz1j5LJmTfuHhEkXzYrLRSXuCLEVJL
MNXkBgLh2JntfF+HN7rw2Ynie/TPBLxqwysRv2DJ+Lwmx3Gubp4ZSuKxp1Y4tajT
5PvT6n2O6m233c9akGTKF5aByubN1fIki+hgAlVwt5JmTIiB9ouHWUStcynSpwWK
pP9e/PFJkyoQ/ucg2qLaXDgSh7VN10tPOTqMLDLx+FNqkXPQT6zuQBPcuxmi1sJT
TukuuJGFQjLZ/K/BSmLn0iXk7I+yKDGaVcmJHZNhs+zjgwdmOPTzIBMkKdyZX0Sg
xyTZDaWIhjeVPAG3OXNCjL2MXONSh8jCyzBXR/yy+hbawb1Z4kjgC1JeozdMJtQ1
+M+ZuaEwtWV4mYFlQRom5E6FOOBVCFrMtR/LlKp0uBQwaIFG7/lwaRapFa2vywFU
ufCDdD92B62JkAz5TK7DPqINqu5iFtQQhQSKNrDj8z3TH+0cRFPP/tRKviiQtvyK
skPBfWIm5vwkVwltp31I6RhgchF/jNVjvywJCw8acl+bOk+34gVrSRkdC3H8wcaj
j8Zz1i3LlWk4bPLmwpEs66FpLaiLb38HWIhGPTwVpedaD8k0YlZdM4v3lA5WmKRy
1oGZG98ozSgbNMlGirNwQw218P/mSzKdixCPJ8HRkSrSw4TV2Gzzj44FSU5Ia4Ch
l2Rpf+azqNJwpeefBvBv16bsTMPRTWKIkADBQu5rxG/Wm46gsLkauKhc3v5wguuo
MGJP82RcQqfsFMFOYm3kE/MK3Nuy/KA6KPkrih/W7BMwE6r6I2ZhrMI3GAwv+uMU
mfUoG67qMgKLFnDsx1RnsKecS2piw2XUsGxt1Wf2GqPWWq8R2nBEPgGQsBQaqQT+
9p+9B3TFIX2um21vuAyUq5nYFrBt82FiRyTFYuan3aYM8llk3Cy/bJ7B0psMbbDn
IYjBwmo+DM8cBTjwGiEKnFEBSSBuBuCrbAVWLUUliZ4l4K0tF62zokhBbA+8VY2R
cxip0OXghfEEHYCnQBcqzBhAbsmhJjgwk3z8VsY2ZnAHjmzUikVaumF4iCSGKERC
/duncNRYbnjo3wybrUH3370jA5kEON/ZFEP9nxVXMmpmwZ35CbLc/lQhhDixKe6s
YvtUIOlRQ7GCZnLgmukJREg/MHu3JIX//UgUOxTtTNM/Sr6gNjfwtYHQCRltcwrj
BJoQEfWSrXVTB8Lfc4wjmdRjyzoR9FSDOUISVzfj019B4Thlr244AMIHjfTbqWLB
jn0TMLDanJCay9fBRyrJhLBZmqOcrhWe6nHCD7+rZkNJHXhaw5BAULJw109bjczm
YRn7l1jA/vA6I+SPXvQApzOFLE0msAd5Ld93FPzPgz5J59dZTVnBwVQo/5rUFbq2
03TsUrEg2fZJoFJV8ZMXaYxQKUp71+cI+tI6Oc9dkzVuTWDmrR25HxQOWHd6M/ki
7AVcWRZaSchMeLsTtDNV3CIt/FnaAWjZSsqURa10IS2F3/NIc8Z18h+M8YR1ON2m
r8fctJAC+5BrUtAgDYg7yK035z6MM9aDLjX1PF+80otayAKU5ybRkauopdbFeNvY
Nfal9Mbd1XR6tbKNxIuakkujGwgkHlcE/1YTy601tyq/p7R+A14vpGnmebbWRFEe
UriCwbI/Hv24abNic9zJwLM1eqOh4KokKzg1abxPYfhI2d3voKEbL8VTTa7zMF4u
hEgR7SRuXP41fu+rHLmDnTUAmFq8jGO55Ijr+TDkVzIK4A4/7+3AtbfTZoPJMhl+
t7nGyfvguYT1Nqc3A+RsXM+bsFsdUlpobsq6iSLFeBRn5zyyHsSQYTFLjvULWV9i
0z8h9228lTy6y+t7WIdjk6kBzGrJdqSxPKeEb1Wuj+ICMjctFvnxRqnXPn0G7SOb
MvqAnwTJy7fyZhQpKKU42UOefkBIhIqIvixjtYPJ8aQlxMMcxOmmF20s+e+4yrP3
lLkaiSiTeJHQx0OGV9Bgpfw9jEfakf+6jbzuqI5+MRW7ssQFCkCCW81nrEEJmx7t
ckxpnZZJPKQjPtCK2MtxtyvHN+hfZvhljIvvsLLAWj5lI0/RcfLp5Egjf6Om2HVP
r1HU79gXT5UE55YyjGZUUlDQvpDX3YTM/1bR5IzqbjnSBoC0WUdIgFCD7lNMHIPt
rGnBuwCN5q4YK7qshG04uuUlsho0B4cs/KLPmnJDcQKO8itGz5Ss5s66BT/QOv/3
f6PMj3xMLScHEWB/rxHvgYdjGqKBe5zA5P36buwGZx7sLCoGckMNPFErzdKFyDPB
8QyggCdXdfvnOJB9r9Ft62JvCjGcBgLFLQ8ONJfpBW2NMFl8KdHetD7lbt2Vmrdt
ZmHjvmIVdx9SBaiHisETDkMXo4bgETeI0HBZ78LVrTy2JNdcJCgBFvk8f5niLVHD
HtvlMH/e7TKWMZ+AQvU8HCXpeyLinPeSRtnM09aoW3LVz+VaUAnZ9+ZaCdJJRgqi
qnqvnkPLRbuawfIKrp44m6ELtL8gA/JTtrfo/OUgu2klU294xYfMtT02LOQcRYD+
NJN2Kz35MEOzkQ5Il5xVdI45r4DADIjQRyESOnjOr7CZwX/Td0Ew0ySNWrWpsb8R
s8vs4UggbK1X9el2InvAcwj7tK00e+w63b/xKCFO56glbmq3zWunnvO2ipzQ7VDQ
iXsG9MQTC6/eryLfVTCvkPHRCvfK8TwMAoUXK8CLpUNzp+N+ivADYKReIIELEeGQ
r0yKUgUx04x0zSfxjNDSFkYAOZGB2vd059AVsFHhKcUBsrKBFUnFsa8jGuf6bmxg
C0YR4CclkK/SEWoXK1aKYg+qrqR2TonF9c2Ba3RXn3MxEwKLJq7tmNfb09qlWa0I
SnnyAEaAbyJS5ylGozLb6fhnfJNyjMB/UI1qipUSvZVxt1fXgeYQ3BgOtGUnX5ib
9LxbQctOZEXtnh3Qn5OJCfbDeDshTfyFTQVuNWR7eCWH6oxhEtcOXFFd5LUqlpPr
maUiXWM4OxaBwf+6RpJsJaBAEbKeNiBVwmNO+cKfGohqYvu7NvrDOSFrdU0Qfft4
GkLy6imkbRcU/sIm/VhG3N09U2hmOlpEXJ7obMMSa7pF2yLIz6e+5vUUplKSOb5w
kFjqKkekjI1aZ66lfGq0JqUEFFXCAduH2uG3dacCzN6eQZwSNWoF9wdq3Zlf/di3
tY1DNh9nXxX+/CPAnzk72q4sKq8RSkS83vrPa6GwpLaCSo8R1Nphtc8K6mYFz5eQ
85vB2F7o1PXqs7QgHo0OsZI4Da3T9mStCyXxp1ZiXFcMUr5CX5IqBBk1WhdzOnMa
s5Hl4t4qFUN9+p9VnszTQsM1vfvkHjDNYa5pCsN18tfrVKPCWKn9jlrTDxO3si40
CyOSEYeUDVLRuYCYpkhRh2cJW+ZaV+iXSLpm/WfhYn4+kYBox0O1kN25wpkcZ5nt
iK5wMMe8X6oFb63CafE0pBb1GPUmhH0ihd8SApAleasel+M11sFrVrqjU1upzj1q
Ul3ziN2wNdQvjbK3SEsNSJez4cCMHxIPh71cHPvpik9AfeEVQ9HJMYO3KKa7fJr1
53NEzb3COax9PcpYApepmCD2CDP7tYUMJzR/jGXeK16nBaldePemti18VaeDnWhD
JonDza569LBVjIaUzQJ/FgQ6AIv4t2CD7wHgYTixzJVVBLp+BiNoeoGSqPkOHqi9
bNnaLkNp4oda8DODOBJAaJQP/x5Y7EYGDE+l2GZBduq3Lbv+PLGRQooeNlgxMDBe
HHNPQQtBQqWrqHcy2KXMK2JkGcvY/h97M5xVgeZK91BxTJ4HdK5NZWWKwOQ4lIFk
7ETOnZ3a4k2VNO5lL/+p8592Fi2WQi29J5DOQoDmCnFRb+tD/w3dGsj50/j/moNw
PIePcRmkQi4/U3fffCo/qKyUr9VGwgJhjRVfa02R9UmIbvTbwKK7fqH8a+l6Ns8+
zthJioAM7Efl22sY+ci82s5lO/oHlEbeiFg4ge3rWot1sN5TnpQ5sK12j06vZaPe
yPcgNQVURJfREHIEubOH5TQyCBSu9tdUVyOQWVttXR3ZkW4IOWEBKsQRirOnqvjq
32HXD8jurjlSRVvj6w5b2kYxV8G0Hhdp1ki6Md0s0q+mT7k0ptA6lYfXGUBOkd3Y
ewqag9MUXfzQDJoSLGYxRfFvt2vFUEDKe6BRG/clMXLyqkIfurjYkkJ73xPcKqK4
cx6NppjeHz5g2GLiN8tMHRJjXGaWasO5Id0/YRTuFU+bHzSSkoIfU+bgx+7ke8GZ
y/7/MnbItczFp6wjMLB9+5eJ7sX1j7AjVTxOHOJ50hx3MX/cKAiXv4ISNMhwMpPO
fBtAGZHA9cxhHFccq7A4f918fnQNu2TvhDA8rH/dt6AtRBNNcaAHPTFMJU2gYTQP
F9XeCjEdY4ymc2WQttUOQM+45G2aDM8o/n68qtSv7Q7QINYegGmxVdKongve1kaw
4MNpMyZ7ldYPTQOGq4/U88ANRnsBIq/ifo68rmNfhqjcgLakPEXK3K6pRLf325YR
RE5lwAuOkD/8/+XB1e5o8pR1kE3mMDsyBcov8D9cWqaMOhZOJk1byDOlKtMm+YYR
tnl5+me0hgNqEIsLNOj+JPjjsNTyuecnmxtUXLZJEvnCerAQTE8ZPSwDe12o07x2
NoZhFxIeXB2dc3C7RR+ktNR9qasu/FLb3iyUK/BOObLTvafS+yOnTIGpfMuvXo5b
npWuut0+K1hpC1AksovhMmNTo+sV83Awl5ogz59U4B72OcqHpg1bGbYK6efVXE0y
ncqzDUqP8fruBLylisVpZ9QwuvC31XkjnK+eA+Se9zhzeVfuabhzErdfGSOrWAwx
gYX3D+yq7y92ImuAXmvQVY7++MRNE+V4h/a9VkWf8txfwC3AF7r2CD3mHTzib+oI
bd4nmdf7ZMNxV1e2fpn8iW8SWqWELW1A19ZZXyfzDSd+64rYsAxWsBNtzglqg3SP
EmPPrmwl6AAbjvfn1kdNJl8xv9/P/49wwb78hgHxxJbxGRtmI8rjpbtkzpLXXjQk
31Wz3zO8YS3o06iS9EWbnEimBwyzfElJLXrEQSsw0eKVAsqeZu47zXFqbHdkg0mo
VeHMUIbKI5nAxb3Kg4YWnAdgtnoWRvtOIPbddBPP17hXLZ8E9GwAMw4O1QMNgSzN
3v+Q7vyMo6kfm3J7d4teG9fZ1FYE5p2j6ZNZx7aQ2BL6DyZmB2Be7nTifDsryElx
Nau1sJHvI/0ep+a/Vbagtvm8Iw+F7JNXkrmkYimDlyzXmGuWZ5h7z1Sg/v27gW8O
MVS0hQPVE97BpXTd9NUzko8Wyy4IQA5kakfgAW2bnYTYmBhyqPLZFO8Cjr+feDpR
sK/G2Kb4f9q8ycEaJ/lefTMLdde2USMsTgTkx18tVCxiQIEWfvNiaui7SjuPGbuU
ZqDqUWz0o+eUkyNf8E/3sBHVyfeDQ+1qJfiIDB2cI/6tyyHf8Zi6j8wWWLWz3qB0
s+T/P5VWs8ZCxhqNUnyVihJQjr57LqBIrB9WDWSN1/589ebwo6Xb9f3FnuUa1xwZ
KbN0QI1w7WJ9NNqzkz95iJG6Oc5WdqGBGsYlbhxVaD+9BdsYck5is1+8dnQtSt35
b7V+p4SZ7AEeXPAXi4MD+oqtsqeSOAw/21SAhntfaHanZ8jzaHJxoq9rix9JOknp
VSuV+9A3IJAb2giGfewGJTolGwp3u+T/4TJ8j+3/8W7OQqqKY1yA/p7gt4gL/ZLu
bdqJD2hybDQUEiMPOXG1cHnk0HEAobCE1mkoSsrFokBoQeoY8SMs9/nHXyOLkAgt
P8y4XwNmkhmWDWWIWoQz6nfKMKmwLWigVSCzTbNXF5PvhCukfkiS3nedUdmvvGPA
mIxI/7MEq+KgWGo7tXhZYHPEJ8rDXxL0yE8dPTcA0ewn36wD8NYRRbtU+VwHlOdE
CEa/kLpyk2DFgOQLrrR03Y0YlzJ7OxjuTiHqGKJkDVZw+MC1zsnQIyuy6KBPesrC
MZ+0tj/w+FxHmEU2pC1xd3n3l/NIl4TYNaEXDjKuqAaq6W5bZScz7HfrHFIsSVA+
PFlC1DMqiw02WeRZKv0c8FGmGe0Nph/zEoMoSeqCHBNjICfV4jJu/fNXHaWUuVSS
tAc5zKo5Bakm/fYKD52gf8NPXNH69SQPKD/JZhth8s9hiCA/+jkzBXxpvGS3sOH6
n3biOCBr9Rly5TLgqVVxwxLwCOtHr7hjVB5luWrj+G+f6dpB8IGZ6hjY7SORbkw4
PedqHHyoVJIYpxRun2Nu7d+DWjq6rhVjCBqdw4kytGIe3+dSaFCJ3fWiW0yuXCQr
QZ1FS8vh/AcFGWFI77Wvv08Wp+4FF9z53yVOdm1tleU/E2yFyQy9OBSVonePxH11
+Rjxf7HHWTDmN7SDf096UAVbBTIFmLVW8m1QH3CHs8ohre1axz100qas6F9njDe9
tqorIdeg1A2cKl+vbiFNRmyU7f5cuLY74lDaSic1kI9Mfk1jjVcJLhjs8npnSmPe
hAk++2vdWa0nfi3+rnC2r8Nm2Ab+XqXgSRpZzWuUs5ZLl3vRpOc/GPJ8EzzSDLi4
7lTaAw34cQiK3TqAEAZKpWsZTBzTJv0QBssWEyV+qnuoQckexSBYtoriBxhGIB96
mAfKwLgPJFZDr2nkMAfpUxw4G8IbR1Oh6aPeBRzBVSZ7s42sDAmgw9k4APmJc7h1
b/FYEN33aG7WacWuU14VRV+bhz/nWSqYNmuw+mRVkUEDYq/xkpuA02sdAtOgXgZy
7nm56lJSojLhpUirlD6Fca6x9gVNjrjAI+GdI1B1NIxTHQNp/t0dPez+NtyTKHX6
cmNHQ4GDelc0z/QP0vgHyZaUQ6K21AQZK+sM/ORFksoddsqP53mTotrTJ3vVEja9
3x6JA/Bws3syIdPVhNohLWPh7iwtOC9UP44FL/WY3K4k/jxxsg1wFCmF2YsEptRr
jEL4tFVJFjb8TfXDNvZQDQvLAZFBGQk7T6Mx17Kdu2chyRjKiZiPfD1eHSb0KgaW
qpgFQ83LT7I6O0TjFj1JeMLrruaoZytbsJIdSbcybIfNzpzw+yDqp/M4U4vVgJM/
xYFVikG32yQJ4ZIk9X97F8idIZfRljt4JUuHgg9ZYmQxNhZe5HclMGJnqDrouRbt
8YMvSqP30hdl8BV6Un7ecWmPwN4l/6M6cn9VO9ZwwFCbhqmtlTmcG8KbSLW/FfWU
fwr7mlho0sJ7G30fjXWnVBVBhKyc0sZtqo4Adj06Oq9+Vv/1owJKWAfl7T0bXbgT
PMcfGdCtVuMp31R1LIjNziQybjZTXPfdNsE6/9oQVneXiRmt9xV2Ncq+PcXBzp/R
Qjo3PMOyID29DFV2lSMRcsi3TkJVuWN1RnAd1VAzSG9WxFmfxEfrXo1x2k5fFajV
efBpfkn8S+bnkkUUaAHFWQLPVMS9Rhz+E7FeEz6KUmxhWVeF+r9bRlfUYAfjzNJu
k8ZMipOVyS/qHdO3kanoyPxFw0aoDzv2GBFDXP7nf6Tj1Yy0NjhP1yr+tfe1ID9F
TWN/xpkegzwWhVj/qgJgMFJX900lwVmf+P9+sPK8iLWakuIvgXSwfWpjlgvow4/X
bkKFP8kcMNzqqoJIERElXO6lis47H3wREZdmGBWr+Z/vrpYv0pnBKM27XGs3UuhA
w93uMpNOM1w2aUA0A8PGROEagm+xCyNxxuCjwOwNYXuVpSKUmlKrAeE/EZk3uoXO
+tS42zuQeDz+wV6hJJS9yL7N3O7P0+SEIUFZfyQjKn9Kz5Lbm7Or5kRGARJq6d1a
WSjE/d26COPJlILtlRFhV8qOwViHsigWhfX6drPCpankvoFPiq96029SEuljOA4o
pVMRmEUhwC52w1fk6yJmpd6H/CgwW8kMikj8/yg96r3epDbZ7x57jKPnH3wJoaXq
1Xr7PnMTsJCJC006Du6xjLAt/O2hRRuJQWE6e9o+Z4cgQgjiDNyeZsM6au52d7oJ
IHBMn6tAOfyLAaHF+7ULwNGH55R0nA27H58AegqW18Q9h1LP4JgAyp5I3w8ke9is
3u/UATHAeZsdAKNssNX3+M5M0AU/uGs1b/UenqlGEMFYy++fpie/QRp02EsKVoLV
+bZJJf/XVr47oHdhF+L2y/wrYraneSTQ+ehiaLt5NNxrJJ1sotGHvQEDBZwmnumP
U/cuVJuiuGvpw4Tf8aj1ncNnHcsxT+VW082msIhReho0zD8O6P2J8HYF22g/Dz3x
NbqTM86ix0dqXuUwVqP2/VYthMEepmFtClb0jWh3+pIP1wTavCmUZQ8HoWDrdaNr
gDJveeT9iKibJjBFyVg2IaZ020VoToRk4o7EeGiYq+J5a97jAKqGzJh2Vkaa48XW
ljsL4M6kVci2vHtEY0tTarm5QLqKpiuQcKff+/8jBjCsWAT1bSJYBvOkhFmHUaSj
burOKPHaIshwiYf5lI/fRoyGwDczSWdYQDd93rhn410gJS7p//kLoTM6LtmSqpXk
qqnhjVdkIb3OYBgIt9kg/3afZNMguQwXlyRajjy2llYVTHOVhQRHK5YjA/BAcFBU
rWQr6hiizqEjzd2+s6ij65HuXtTEOQwhKaJOm9l0OyDDw6tEtSFxkK0AxuqfvFMI
O9jXuEENCtBuCmt/28Kzd+oH8BPvZnpZf82P58c7znrEYy0Tf7ly+m27oplSHL9I
O9kIYEHCYcIlvz6bQ+4n15s0lw2ZVx9DJ5QSFS+Lphs7Crv5mbqX43Mdfbo2D7G1
udYHH13AFr9dxAdl3va/gxNrBiYFnx1wfsgn5oa9WAXnfr4EXOBA87FS4qPfpbgX
xCNfBDtQ7PEr3iaK050ivKXkXx9+CmzhVfNstqQwsfjUQ1eT2ei0kqX04BzPLAwE
Uuj8ToyBm2wuepkH3oRrmw/AGglV7S8ZH/Q5t2cMkvAtLll9gyz9QDBeNHxDbM2S
tCwIju6iSgMyuKRnAg+1Ck+PQl89Rjv94C17r6rVVl8HPEYCON0StRzKuGckhfgf
7orzGTJxBiB8kR99vP+A4qBxEZ+2SkZAqXtgfgJehKHoWzTA5ee3tlSm+jqZZNgD
EyAYi4Nvz8oOemuGxBpuWxaD55gUXk5Rmw+YzMgs7ZWHt8nYp/NZBJlTocLfxZdA
RfIe+MGgACiGlTnFbffyYUR8dwfZRPdfG0Ne/8GC6ymVybL0wceIOZGnhsnUI/01
etnnjZMbMrxJptgTwfSNl9pLOeiJQlsuXmpCgh77mxEPV3KWnHqu3QhKCyGE5IEx
2aBD3o6MfQWwTz9LkRCT07vyxVhj3sJcFxDWrLj1B94bWM04ODSG1c+ZVHaPXjYr
oINl7OCWyrVCBAVdj7ZMyWrytTMZ0ROIPHwYQhQ3Xf00TlAm1V9QzRvP8v4fr9xl
Ds7CifmaJgA69X671JOiDaBntuY43cphCWmYjLRVmD6H+JCYmYjoBvubNDmVPLje
TuxYzq8HuFGWw9d0ESKwUzBwWXzGyhni0nSa4UYfzDb2/vfosjDjr663KWyg29TL
MP3aomWUzD+GhY8WLMj7EyW3aH8USUAph6a/FDSicz1KiuxzbO6y4QBrk8ypEtxe
EkB/Dgmw9ZuRuAr7scq0eAXgWf1fBO+/IMU6jBQhtkP6OeSiXP0jzAWcj+tKUQwP
4y8QYo3ZaGKbGoWufUzIj/AQWEgbkJmHp7BtpGPVxJ9IuswWp+M0pslgTCVO0Pbl
GiFWPKoz8ZZw5y0nKmjgexRBTGMvQxH8X0BkeyCU5Q7HUCDT/9OQyLtSBsQioAUA
LawWpElbNZQO11L0qeClqKlIzbDqoIukB0c3I5uz5zjkJzp29UNxtrSMiiGh0amk
Nk6US2paAhoUuqsVSgRmIJZUbSakZAvejBofN/00FWMJwMEimK32fr9GzHJ4RMq8
H8sfbZafGSQ/qjEQ7tr/rZbjNPicC5jA4hbGqqPFxRYrqzjYqUq7xebthz09bqAc
BqA7bDTz3+QUMM3sKMS57AAqP1xykScHLbh/LffUkKkS2D6IEKqNRYeUNPzE3EEJ
FYY2s5mjjWJXYXkgD8w1/HEGYHenoOYxGTvd+2XPkRlz4GVi7ZW25Dt/avY12/Kw
xp2s99LKF3lOnlr8QslUvW2aXPv9nyo5s6PA49eAg4oMyIfMaTwDxHoAvsDB7umZ
Bs3QZK/aSY+Tux6t9msW3Zy2u2QKx1k+lU8OBPNoIijY4FSXKvVAeKmzuIUtqjMg
3201IgUpy/1g+0CpAk9oYJWehdkC13Y8p7WWZQ+La43VFFgi7NuuR3kvCxDvnUZl
kI8CsS9XePqbf/ftgg/W0Rkk9Qhi/k29JSM+U35L/B2Ac/l/xg7vgg9oLvlbPR0O
2OUEP8BTgypj1EQ0nYVw35pxFoM/8C/Cw2eW7YBm5HiJU+/YNvUG8tGZ+v3JajSg
uuLLAHkf9I61J5C9m+BvHt150ZDBIk015MkRa3FFSIzH0hQ03XlX27KbreQjzaKf
EBShiy3hOzkG+G6JPV1DVB1WtaOrbhLm2Z0SNjAWlwTiu4M3MFOuFpnjlM9W9SyV
cICj07Stc8A9lhacj2NN488uo7zip3NYdAFjdpbmiu8kc0NrHB1EPYJpuyAE+0VS
vaKUO45wuPTCCBHk+ZkepfiV9yQp8WKv/nMDlY6jD9NJSC3sbDIJYb4Ln3WFLewC
3dbaiObu4a4Dh6kWsooFqw3lAUa7GfK+BrMzNFXTboY3eY6QFaitGCOJwr6lO7tI
6J04DdF/FUSwCW56RAS1h3t5gQUdsqTEVm2oPpQOMTVSscrbHt34CoZS9D6cMYcy
I5tEb2hNIPz2HmSKKbVSVjhLA28wK3nGWNPnb7x/0Cn28Cd9HgabpN7lct3mJpKI
jVVAkfYEr42rNCnFTrIPnt1MSMP5/p66hEZNruevW6puVomB3X7yvzrsNs3B/t7T
PVVMPF/S7A2nGEIzlGY+fwpehP0oAVdTvTLWNbBeVKx9DscE2TvtRjMj+uh8NGNu
mv/jLP9dqUIuzh2RmXfi3k2gqZi6SJSOxju+14iOJrxm7Q0lA8WJ0k2P4mahyqak
HjpBuwuUPk+t37YTLVAXsag5H3C7gglSW7TYANjA1gSVq1O/No6/iKKhv8YgjmoJ
HAVu7LD8azSu0jGVy3zYm5hxyFKuqGeM29lZPvVnNlEE2NAafcgAlks68kBk7rOo
SFCh7VOHEZPZNCqw5zI5lGSfGbFuhjafjz6ONwdzcKfjthoBgKbLNdq2jfAJng1T
EVmiOPynv2Qv8vpFuB/c8WzfF9bi0QNIQviSQc+3+vuwsYSdDQKaUNSqVRwezJ5m
vbqevwen5EAyJjjfh0GuRBeuA3YAHYSstJtltNIRojUgZxUoXEWA6qHOkI4nwghu
FNE9SOUF/0rQIXbutuKen+tYo5+ZfJnFtvuZ+vHh5eHM46jQoW1yHBwTTnG5Q1FZ
PyEZNOgbOcfjqQyt7jHScBl5DUKEocpTu2EmyDhfxtTCnCzhpBqc0xV6xBEBj+It
H57/B4xvoreJTU++xj3s5PdKOTZ0LzJmXMvuXsXFEiO2e8+1NATfcbihxsctLBss
5A43HXfRCWRcB17jolS8o1urB6Rz2nKKwKboMg6iWSBT8vID52iJ/YdIlUGtnR0O
/2h/7RNKEpDGeq/H+tmv024svlbzWJwtxheNL152ozEZAZMcV+OCUCRb2+Qt2gD1
GIW8s0MG8TtfETQM8Vr/zncu9RN876xc8CfGPnF57v//1F+63IP8bZzh+T8EML6O
pzhP2IuB1RreqJJY4fnWYkEMkVALxdp9bV6IXvjW5vXSDcgsBK/dW6/rrVsRkBrg
wFDs8LmCimtHqHn7D8wFFiuWyWHgmA5QfUWQn0ZDz6DIepi/QKKix2ph0SkeHdDv
MWaoK6HozQ2fu64lCE5vJ5GjSC4tm2dcDd0AQGoLovBAnhMcQyLyrnSPVSrg7+MP
3TrIelDQDcpIhZ70cTy/P2JDOlii44WSbJsLnK7KXydkmVphIhU8OxiahV7/coUX
r80kwAeJPXsGVsj5r7nBytu5U7AlDPEeIcLdqCrdHFKuHOxwZ6RtCR9qqfP8Joon
CsgI9GxaJlmmLIzYYAiDbiW9FZJhdN4DqzjP1C6OAVDoN3RZftLnquDNAhPooSC7
36QKxIuMNIxgelXlnZY+lju/RGLKhAlWmfM9er+tOkfXhFQ6vXdISEm090lrD/mM
KalzuQ119PTUXKoJF7p+EbALoRDh8JP1yQHRNRHAcEV3lPFg/Xe8hBjB+JvFyC3d
QRFR3EddQ0aMchzt3irEPUAIN9wl1VNjIdP2TfibyGxhECKVwkoJH0s0MgC0d6K5
G5676K6j4aDGQZbJKLxg+a5/Dn9nXWV2wzqJxNg/qYMGdCz2i/jb86dcfUJFJ8pL
ABFry8XTEbur/qtjsISTpY6b2ZDrhZEHAlxwonHWL2sAl4YTbQ1Nf5wCPYeTZcrW
xW+Jl3BjonD2ZZ6+6R+YKL8H2oa+IQGUdHv2SWWbSrwGT8cjnEAz/0SEUxF+53yW
u2n1LdqZE/qTXBLHuQd3a4FNfEu5hgqQuO2EP+h0KPnxl9DK+N15ulRxcisuaYq/
GETVhQsbXQ4MQDNQWOHu/r7suZgNSVWcJZMe8nquTWiEs7fikB1XfK2/0z5I4oPK
Q1jmIgl3Sp8z3nIhNX+JCjxlz4aP8DyKzvppyX9KONnRa/1KuSpP1vEVBP9W4jMh
LZu7dcS7fJ+TX+cWQok+7EWXMsdYY1HlS28hpfbIdwfnQTfEjB63DDVWL0LTtvPS
hdr7nBbHmgzEBqemMjOWBJa1nwzo3eg8cnKbt7KUtfBbTkmRWjcOHZ63lFNG47Ji
wwJCdXGUWNgCI/byFFpKDNp2joql4BcaQKnQLw+Dk76uJkTvZlgbL7Kej7WDvlA+
Kb+XOZ8OpXHPInFJWXGTR2qmER4AfM6mMs5GD8PsVpCdkhzzdfymPGZyOEp+H4ER
RTBvmFyZiBznh3Krj0O73eCJKi1md5nalyuiQhkSSEzb4ce2ar+9n4dse4wnKwKq
I/zqMipa+lV2B6OMvSELa2P2ENJwD+M1qwnoPuGzZsGAj30yE5LukJ7MyiNIWQRg
HHcDRiQuCxHPqH6NV9SEkfPJiMS8AbhAsejYIZddscHoF0QvJdF9bKdye/Kqb9qP
EgAWQlgQfHrA2KR6yxDkXoiye8ji2WmPPsTrKPG2YE7EIGrDaAWBc87ahxtbiaCz
ebyXW7KZWG/fn77ssWZxOjW1e8A0sC7UA+b7El5dMJQk95UixvHrj/V1y2jtRA0h
h/dXPRnPd+Tv/bdU+SzsUwt4j9EA40hPMLlhRjEsn+TlxK+n2Q2CXo7mSKYiDH1r
j0IVdovUrQpVxOIUS+M2jmrrvmmWD1HHKIwBkYW4bllwvc5x7M07h9QeRbsRhl+5
zh9tbtdZjeomHpCiTJdYjWpoc5Qwj0ponHinz445NsL3FFzsxwYmYAzk0rl2q4MN
u3M3NVwl/agm+lhMGZQLzGvnY6Mn7aUj1vqapkdqIj6ItwDKPlklIk79NFD8AI9V
hhn5yDDsQD2E3PZBNdGlg10O6kgk4qJxXfsqPvLN882XVZLPrav/PXLpJ9+QnsvA
nTfClNJ90ygTcW/NRFgCSdEOGwRbT8I+iDD0tivNrhFTzKKS5c4s6I0pqqDXpCBv
l+JVhOhSUBKb26Urg0MoHg1zTPSYBnFCTncmOHZq0MUCbDytLgFzWm3AyxQflruw
s2yLcXpfwB2P/Jn2r5tR5mQPRlUxqeDMu4Af1poPi5hVDA9TNzD+TN0/Dc+vasoA
Xan2RsESknRJTMpC9MZA/XaeZJiNWRbjG5wwg8Fk5KYyoAo1oEvq7qOuTZuVC8aS
AjQu6FtL+99B641S0W1sYUYrkTLJ/JBS1fIeALUdBAJwdpppQr30ofWCB56kzbaZ
WkEQwXDKo/Xl51FUUc64ek3ruwbpEgSOkpxvFltoIqRTtN1iqpou4x9tMCCLFTnj
Pr53uBhKM9+174RwpIT/2otK8+AaNJ6fi0poMBTKf7sETjDDiTDh7W39goOUM+Nf
evhohHAxydd7eJp7d+nCPq+DO4iVBxOKsD2jZ/a26VjNun/2T69NZlSnG/RhiXEz
slt72Uwof0BzfmV+PekqZ67Y0Jb8/t1qCYWf4viQmj6VAjE0TYct7yv/2mAlmH3U
gOvro62V/pIUZ8VlRxWGD0PMwsPI1T0qfseIpFfSVbkiekrs6yoSRkakau+fB/IL
cdydviuVZqMcHUL95yxk1ExTaEra55a2/1PftizL8Nc7FSmFPXJMJVz8uOp5izXW
wo7iwE24hbWHFFrb56jnvE8A1a+lopH1V7etxqhtgvHaPhDK6stz8H/VLNagvKsa
LF4dY50Kbzj0CpVuybw7sSZ/RqLlfXR1vP3XCCDpKIfXjVPxQduTmxVwENOjuCbt
9/R+ZnFiTe7WuP7H0LZLioDaOxfBOs4C7AH3Vdq2n5zZpS/14hsZo2Yk+WVrWN0X
7Oe/nbRMJ0TmHaNqACFpesqEUk6zFcUyI3tLC18Soepu5KbftYMsNWOryEzeDdxs
mt3HQNmu6lBpe94d+gGoC0tw2S2oik+YWTMAE21mA/QhZX6jsnKZtthmq2o2Rggg
grVmQQCZ/Tu76eMq5t5phZmmWpFyQTfjfdb8iOy5gGRHxnqDNXaUkNnAsQs88XqC
pIU0AttG6pX0OzEMQXDxaMzYrmvbZBUR3NcZsgYZF4hQP+sxSfvqxPRXtIXzZx8Q
hs9w1XXdcnLjXdivqUsqL+MixMhnWnqZaTlHMel20pKMqcU6iaaYYt05AqnShtWT
77MSkhj97x4GYdd76CWjVjHE9resI010xbA16QL0TBqz1fOn36dYV8kqcr8iRiz6
/cXtL9mHZRQYES35vl1XR63XL1B87tlIl9XIW1KBYZRxB7f0oy/ou48lvYuT5Pc/
0AiU9NyHn9QCRTh6mAdhCtAFUtMyOxToqLsqvNZZ9gDFu3E2ZW+0mfzXiO8vA/1e
hXcyqsZ4+DC9gQ90jLkwUQ1nDAWplp4OFoYxoxaAKqR0KDlVOzKbzojho/VMBXiL
oWxwZpo1Vczif4+ezz+XXBUa+/LHyjWAZ4biQmQI8Bn8lhBbm/vMiqOTAZR01xWj
ndYykhRwUDEO40uVVhq11iraBR8H8j+wUI4wj8W4sqRuucDLYRhVkD31em0Gcrg9
7sdyygbaQ5F6xCtyoSUxHRA5JdZLFS4255tOq2Z/2rulYDEx6/y4Agu2ycKnVGg3
wTdEHcn1gxQE/dK9p5MtuiNJ5tilSKcoVajcYThLz7mda/ZsdXWVsq7aSxCsdl3Z
tMJqT1jHkIGCW0BZ/Hd+mZJSa4XX1fDqVtmkmv4idyqNQnUD1zZYpRM1xAWXFiqS
uIZHHaE/AGkT7sFCwGePNRQjr3Hwp4rlunSUMFu9cZvZ4Ux2IUOPz2kcfdZwz0Ez
DASmQUKm2gsX5hXr5mHOX+Sltg/KcOT+cFsSIvxXWexE5jODb0/QSNv5k/UMUrJS
UWhS3t3T6nukRtlB13byu9EaolI+s7i/5JaWtt4FoPAj2N7H/Sa41waGXTcLJSyN
T+M6JJIDlmW9Fyd/YMI2d2nhYNdfk/1242qJBrC5ENWFsHs/DuDmehtF7vpxe1Ju
8z1aXYKGd9vKw7ZeXEaUZ4zSX9v0OIDFHmXZT5WOQx8hCRbPj6VN3TjOr7HHWVNv
xc5MaWIGBv3hlBi2jqeTnutmYX0FQIpqE7adNBlKJTq8lnm55ZIJturhWHQyhbas
bCU0R98f/OYVqNaNl37wl/yZO14H149DJRnsN3Mt/z1j63EfSQVLYoid2s8xYqOe
8IySyFw4dtatM0wp8gkF0h0Zx8/0cxKeNKniUHIeZS3JjKAQcDJLctW0ggFCSDCx
nK1n4BfsAK+Lj4FAgltqrOVUP7Drl7OeQBmPWE0N2Vt/wfUCJxy0gLj/kLtS52M0
3cKReZHixZcOoV/TU12hAayVPsfXR8LMZbPhycZU5S8CvSEXBE30PhIWL6E6rQ7i
Yj4KIOx8C2zTv7cGLpdA037TuvaFGI7IErkYN6BzxO2gBKPV3/78BE3jwbRIedKF
x1S8JXpBv6nMoNCGTeOg4VKzGEEnZLUSn+8K//jScs8cq9Wb7SZhW+fiFE434/VU
4m+Xp3i378Fo3hAmTPh3OzotQR8qwHO68+aeyPCLVru7VyJ/qctWfKUUTnrupVY1
xuEXke1DxLlaDQuTtWEWTcaNpN0Ui0eaVl938pNLyzgho2D/R/vExEVYOoF1lYTY
UZzgqfAOXJ6rdNQ8KVV5tZHbp/4EMY83J2FO8A+DkWp12vY4rPvX11k1TCElJYyO
bkXpSSpu4+UWDfVJ4MlalZcYuAHg4d2YhWVCVpLaxF2aSWufI0eroJ60IwN1Hb7z
VGXLlnngENpnZPzfBw29Efpq4QgX3RtlxwXQWRz/vDo1NMtB0bUsXVJkrQ2e64yO
6xwucyyL+QIFFGLQOgJ6LcHCXsq3ycYzPJSLKDj1AqEjFRjK0BXUzP/u7z6G1fqv
w86eSrjzRoq0Rm2MmFfHWG1A0UB0X1Zi0t9aqLOB66VT8EsSJLhq8HUEW9pV51Ag
ZmeohpcVEcRXVOIXcO/K/c7qpXwiWUt4whNa+1XwrkcrGBzIMJyP5tASdj1a29Fd
5jajnxlRjy1GrVwHRbYfJJMp9ApBawTbxnA5c7HRO/8llvL/oHp04cuG37JR9i4F
5kQezp6Sp39MHTM+c6N6Zno0Y61pXqVQjsaPtEYiufPmPn1s1u9guF82mpFtVl1g
jQfYTqq2HYBN80S0g0JMeP8lqOrgXsbCTb9xYXU1Vneo6Q5nZoTtqdsUJPeleW0V
MTUal1Ka9fcM4Q8qFHcIispyoY44blIoL76jki3O+kuV/JtOckOffd4z63CGTH6D
AhaoQyFnyn6sw9jK2IDbKlYwuOnkbOGfci5UhvliOH/Lr641AJKbnpEDN5uDDcJV
UePWAMIk3+WlLBPIB6FX/phlNWi44kL7nCeVb6rjFx9yNVWwzJniiLYQAYASRv4e
jmVVynTlrumthXxXTwtdnMzw3roUCLgcuctm+Pnf9JX37i5RMvDH0u9omZDXBOOK
mBUErIJPRWQqigUXe9NDf2E/agkFgEyQjNtZB8gkICCmnjyjg3AphpszYeD7zZZ7
OfSFhmbzpkAuOA7qmxbJBK5RYkz8O6XWxOzQux80FiMihBia5YgSt9SeYHPYdcRW
rWbfKmCRGG/Z9Qa1pCptDOU8kcn2mcQJi98HxIE7CfpcZwj6fRg6p5TzryzbFZ51
l7EBmMO+i7yOZIUb6zmI1BvmIEnKkztQcJJ5Q/KQgJIn8IBe0ukkO13F6l3LuLja
nSYw7UGQehrkmY2gntmMNwhgREZ23U0qGhmXdSwQcQQ/Zf3Jco4QrdVJguEQY9ZU
6p4u0JyrmjGpiKCR7428X1+X+Sg4J3YDS8XQJWALjTei6dMcclHDTfDya7br1TMT
rqIY8v/pcMpbEDEDNCdjZ31+bDJ1tRZRqsd+kcUCkMc+nY+ZmT4qtxZYerKcporv
1+Ym9pdKd5Y54AcMzi8vnwLl3toO+kJh9fjRG6syBx5llzOzFqCxSo4jrnHxhdGf
/OgcGtjran27REcBIchLDP7ZCCKfGSdauwyzKijT76KnVW0emR7tWYoTSXuPoyW3
FumNwdhBlYBr3CxNeO0EdcXsydKYTveUwV4hbhpAhfRxoR/zmCXIvFTpuqpX3Re5
Z84ALHbjCuXFf09TFW0LtIlqqY5EhDSsDhEUlrLCD/n7eA6ew+Ho0NojHfIn8LqF
IAq2o1enYEmrIx7sSuEG6EHF0PJ5QhG2OA8Qj9GGC5LFFKXXh6TSplT29I9exKOR
n2f6nVyN5BWKwRG26RLGHavjOqMVFkBD8cz8eNwt25QPArB5dgMDFW+Df9ourHCk
fW0IY9vrgJJ61vhZ6kxgNiDGjc6QWbPqTFx1CkCUaJi9Gw3p1blcn667xPmD89oq
XV9qqmetDGckwBO/tRpiN8FkRgcKwBmrqCAb/6FC4UzoLUZ9Sj9fK77xa+j+xI2M
psviMkTv1zbN7oGMsdedis/ddmGsqLrh712+EVgey/tJiSZxYNnAhgH8TLvJvTBo
Da3VWR8QojXf4PiDijdKGd3I8sX/EpXeul+/OK8eY141ACGxnDJ4fC/dORNucOnd
leLq8fTAAzS8xBwqKCxJFnbdwsfHMYQlXc6Ocgq0WAQPWqt1dq76riwwDMhwX5++
O7D7hlG6Rc6PW0wqp/A1pkzKa7y1WnwbyuJ+HHj1xBIoPndJrVDKyJVoYmaZGmsw
ShYb9gpplCzGEy/42P76GeOtLYrHvHi+0ryhQ7HP/hg6zbtTqXYTNbp97sIdslcC
QGX7ZRjO+ydi43Lh1dUd5qXBIAa61WlMRTpUPJdxBmHM5TgnZZzPMc5cxySoC+xD
ApUgtCZegddGHBXqVMrAMnM0vcPxpbce63rv7k9ySxStgREbp+84tzNQFQ0KFvLo
PC3tCgB8OVp5HUM/WmrQut9j1SHdTpPEFtDI5JMeZZ6R+vs1Dy2kG6J5xOAoDzvp
eFb3+0nkA8hjWSFM/fylSfiui15lGPJqEu4t7twBcPZyIVTW2LeUPuKVMVDH1e/7
ZQsLl+AmwM0bQBYsthq1qKg4f0UY7zpnuPaWmjkR0CO71ggxq1RO6hHEKy14eYRj
Zr35tNLtgUSyNAt0dpsWot4PlKCWw1tOHrmJXSPj8DPlyBd9gg9EksdrZSqqP/6Z
1f1Uyqdwy4H3MGFfD5aF4WeFkPL3CGnOLLKkjZg6TkMReSBKcNkNRJ3p4JH94t/L
N6MyCwfBEq0oXP4kb7DaVX4N0dDe91sqomU3idswrWtLvloFc2StwOl3IUw1GNv2
g7JldGbprjwBAfIZ6QwKhxGT8tbQnQdN6AYFT1CruO+QH148H5CPsR00D0TU5hQ1
lQ5A47OBOfBbFmRMsoNuLnQGgDXqV0/W2KdLjzwZRDi6E1NYww8fIZ9C283yulat
tlmI3BaGPf9tFtgiOAVZHY5/vIoj7AhCZHCE4MZMfJypbAt1JE2ahd8u/LXM3MYV
snJl7MegvfgWMeMKko5c/U7iLRYJDdkwsnMyHi+RrisHb0FoVeIdgo+WISkT36yv
U+CQ0m73qaR8i9qJLQ73d2gi8awBd+sHKP3Ohr1GtWgwPu6+3ZJPTf4b5/e+oszc
xzmsV555LOjyZkEYoe+YQtYFSxbpT1h7p/kwPAwmuhtRJe4A17gXFyP/u9wZrAlv
/8FutCMPMM7cfO45mRCqAG0XHDAnOWBEfRIU1rJkX5f6nbh44N6Vj7ePYqU91CX7
olB4P7JUAB/HWIJD0xETDZBLdN1Rvw69io8ftnYkHYGevhhtXzNhfFa4J/11pX9P
M+oQXjSAgRI1qrx3QtlAph/JnYmlDlGN0BAW6LXC8pjhn/pNo6TcRVG9IRMbBhZq
YQY3eJIwTPF6GNzT3Mh56xsFoYKTJl3ZGeRmDk/EamXYhq/En3LC60SMtjHnNQoF
l76IyjMvqxH1avPSGjuTywz61IMnkwoffEc8lpVnWhDF1Dq6OKr0mmJvj8DzLS5y
wuv2yUtoSBp1Ow/c/P57PmTwlOlzDKdLBiRhgoyDtLNdZopSMwtfrILGg+Oif8Kv
nAdeQWj+cqC1T8I9NRg+BBrxlCa6DxjJFZ3cTHSH9efBZe4gKc2I7zAOfBMIGqEG
FhfR132WLPdId5Z1xsVBNN751yQ7WIYOh+MsGWJUe+MxGSb6BCStHjWvDEQFQ2IN
+9sVvF0+OFE/eg5uP9fvOx1kOkdfkyIjzFBLgFhMaldlxQSoiJX4oxM7b0y3wpNF
c5IEe+PRPErHjiXhcQISDDrlOn7V4XQVqh6jxlJWCgvPBQOR3wPT9zuUcGscrjZv
OkCkGLKKq9/cP9crTO4CcTsD8eFMQ2Yg+tYtIwuGuGAEOlffZICF5a2s41ri2vcE
Dg8+4OmkA5iu2cqsiNcbjfd4qW8+FdpIcMyn7uu4nHBPrQclDaMF2LUeAYhbzI4r
/OVDxHTKwPIWdUv8b2aOnrTpS8sXAuTvM7hyQKg9Mk4rHwDYkePuZkIo+Sw2chEz
9HZr82yDOGG7BJdE9f2iaZPNJ/wRxxyp8GCrhEWAZBi0X7radI6WppIgzuQo72Pv
w8fIPVnIIaAMKUTKkZeCvqgIEBqSvDJKEANLqI2pPmzxgU0ZyF/LCL4Vr9dpFiQs
maZHxKjTkV/Rqop1iGnqvHS64DUE7n/JUABZmJQta6DHTP54zyESwRNtd6exr3TN
do2uHeAz/aYN//GlbPngMIvOaBrB9XLJocSqYiJz3faLfoB0+BRf5fSJXtLTRdqH
/sL08pkiB/LllkiPrS4t+eW97DfYB4nevfz6/qYGCQgG4tE0lH1r4EkgpSLlMOO8
tksc+4hisVMtTywQbtWKwTO6VCUYw4j+rV5VDrvhwqays0FE1ovZgDAO65jtbwGt
U1D+wOfC1yFMWMawyyEun3OR27JyPgkJczPvlixMO+D1Uj91BkhKTTdD5zK0gsiv
JfEuL6/CV+OEQv7eXr2HcvQO55DE+q24r2zv9qkHu2ghuqzKPdImexTd3MQgac0y
DRVyldYdO790zLN9X5FZw16qudZQzNqBD4ExBwvC0PLkjf++9v5X/Rhw8Z9eF4T+
AakHmIbN7zuxaUn5RrGUJqDYJrZksC5P5tgrFifMTQ+Vn8Y87Ei9y3X2lXe6OOS+
7kKOmTwdRI8WHsOs5tE+jjkNxGwbAfxtWtsyQ1y8uQnE93SSo3xkMTQZJHFPdXv0
nlFjTzGAAju/fXJLTw4CVy99q4NR7Wlv61Hhtx1axX2bPJdPX2FoDuw7mlRZwgSZ
rLqz+0GpT2FgAH1Ddc3ptmt7DUpBib4DiP3ICzaJwnD1vt24ZK5p+i6PCuK2ZQIR
1HYC8ecToOfWZocWI6MNIrF9Wvl1MPnJR7Z93nPcrhmskaCYUf74zD0f8ksQ0xag
hc4PE8II1B27O87Pbr7TGDzAf3WCIVRFiTM7EIVuyoVr2wM3rszQiOj2XXy9xu4O
WVZecTXu2NMHNfiAq9qCqBS0aSniMWDWcGlyhocwv86BPMvJSsLi06HBvxSIbmoA
61DfB2/hC+l5QHxw4yQ1glgaNMa1X3+AqFnK7msQYOj/SgBDurVLVJvAddnI45mS
8scarbSQEkQxn1VzfnqFOOq11UM+p9h9Iuf8bdyJYP1c3u9h7jXSOUZL8lfT4z8Q
s7Wn8/vjGJc6mtiOURU7JLx3qO+UAl41gLIosk0Lp3HGMSeJ/28rgkOmdyKH02jV
/Df8qInSknKkjfDj+EywGukk5Y9u+TLTWOHwAJ4VycAEPmwW70aXUSJozZfj3SMq
DeDyTDRU/oPImpAA4TYULLDwPROHTHJHjQK9kM3V5+HRMzw9pHONfp3igixxLGCs
uNEBtMqWx4KdWpFJNw5SZZeHqwo95p+qRgkstUATBE/poaCyB1EedyNNrcI895tv
erCgHgi9vA/+oEI4eO4nuKpzD4888q9p10rhvCa+y2TTRb8B/hUynW9PPp0GsZqo
2Y97fD02lLXRMVxZzVNFroFBzCEz6WZyQeSUUeD2nTxMZxOF5oYTmqMmRyhZ/PkU
J+qLPDbavhe1OfUFdbx2s8xorTtUqPXrroMysSAlabi4pQqH9B+VZfRIu3tPekhy
lofJuVwRCYQTOgbfur2uwDppLogUbqD6puQ9Ii/qXhWGwr3NXw1NP8vHgUObi93U
RbDYJDoUxUfPBtAp4iVpIeDdQW38FvHkKll3MEATTokdI8djcK2DMeGtmrizcrP5
1pAaiOslGJR4HE/Rm1l/0fTGkMmS0+m/Sm9XZoNEaKczqr7bKHQyh6jgz+Q2Y+3i
UrCCgR6ZHJPGPLRDhyYYWkZaoI6Gx6FVT9Ze043txCBt4cD3RTewWwuLH+G/j2nT
JvKdNbpZM1hDi4X/4hWCoZKcRFyDAM3OcDsC+z1JeunDbZIIFZU/giCWFvWE+2zS
QN1y5JqqGBYF8AipU9lBhJdnQcjceARIJKYIXjh5aYH3qNO3OH4b90ohZSpgkIg8
9KFD33uMxbJzekzNgQioETxOuK6nsq1jj8TDv4MB4mvz4CsNgI1qILRQYnUWF/h/
+iI8kX83+KQ2KfD5x7wbLs3b1oSbDCaBPH3f3a77k9a0ckFs0Ox7TTK7AqSrcMI8
PJqQEji1i0AkxtmG6Pl4NIrFxEnFFgGM4qgxzh4SbMKvko3WSShquZS471kxDv4r
f0UGxjYXLEMabGxLZU0OnjBIVV8oWF+8tq8SE+gn3AEtJgZ7R1fwNAotqlgyx13l
Mh/FywCWPdXX6A8/xMZ764BmWnizOCtzZcF5VW6pe3E4zOz2ikvgPtBmnLUHXMuq
T18eWhqhepbecAHG2wCydw5BS/5GhFKMZEkYIWXOI99MAz0/oHmA/KCRJ/RuHQcf
gLn/dcSolEk4Ew+rCYfJ/RCobdsaF4NCfQnDiIKgrQlkg9pa5irIvfQr+1rPhaMX
GkfevDOvuZtknwaCYDpJS0Gl0f1dOZYz/r5rQHpUs5GEM6UNW32nkGEejrRCGi/y
r3lMuEG+nzlW5gL+RwL+/ysGlPvCTK4PdlRndg4GWNw+h71uZc/aKZFRV5MrMfyB
cdqOG5RcLXXPNCe3JIunIk6xPAjLLRcmT3nqIcO9yCo8nd7mWWJgFk5aadgaafKN
R+adzvc4Uk4J2hVa2pG1UwPgzEGJkRmOGtwKgC0UCECHDRcJhObQ8h0bnJNXOnkV
pXlBKCsFdesJDj8sYZsW8vutg2TQQm7uA6BSh8B6quWeSFS4fOUfsmAcdTnOvCn6
VI3FkeqjKQVbpkoOeaQwmzFhfbDYwrWcrfPGR3uCfDMKmVyGVjsYwktJB80Hudzv
DNuxMuepXqpDOcUgnj9kL3SEaARajbObEHzfHkTxo56Gu0saU2YBv7j5Fd4GQoKg
lTZ35FT0zOR6H0oivWZyt41VHsVWOWqu33/m3kPwq3x/68FobEYly8xmt1NoGJb3
/7cqFC9UkxG092CTZE8gdFFvqUC9Ce4cwAEN1pMNJHHIquRz75ZscaKrMbFdNVyu
3vQIWTFhydFROaDhCKNY/2h5zQd7A8CZLoew1q8U2UXqO8V2+v9zJPE/yG8+Qtmo
fyEFMuHRhAjWcKtk78QBS2lp7QYEc/qS23uVsuUnAvHV5tUzU1GDZ4tn0yMUF47F
SQmIwGepbfdaqYTi+YSiEzSQDbBQv0lzDRpJ0pPJNk6t0acLqPXa7CuViCSxPvak
PHD3vU0gq53b+Eh4D4ewRThnqp0P6MuCi9vvwr3q8uWKwGgpuhQAb6zNzJX2kAWe
NlordlX28AhhUnu/yrEM+Z7xKI7wXle51oQOkWQQOSL9R0H4Xrp9n9AKldftdRaK
R5GbSmwxyqp3reHbZoWBQk8TajTewgZPd0BHvahuBhvGgvvO5RZuLTZPNSA0qc0F
z5pobUdPbDVByUYwvjBA7ZVHC+2udeGgOXy7RHB8cFwM+LKFvjbN0/VLkmnwbErQ
dMB1lOeicxZsodFnYOPdK8gOEbsuC1sNiuGKSA1X/qZw1kwSi/slrcX1Lm4dxupY
CnejUaTLDd+IfNUmpKJKab25q/UANMrQ+5YeL54PTh+ZzeDqZSzVW8DzYMmIDbo/
1OtYRzPQMv3I7KWm5v+6TrRTCcZ4ZYS8se7lOCWGIlSZl9F/gHe4akaL+I73rndt
4kXEYRmTbePyKg94qZflyaGBzP5JnJQ4hu7AxLM8kP18TnhHMfI2NXPwmMe6VYeU
4mZggDfSdsfEsj8f3o5JKJO3YRKRebFYLsNLos5ed7IVPKzM+r9BwodMdWqzrQsO
LAZitsM7rv0sAYirb2z4C6UQoKxOfh4N75se5MHsuBIiXb+9TDR2A30TwYIfT1R6
Sw8YhImZ9fINLyl2WcMpCLPsZd/jrwaKYnxa/3mjbPnxJ9cwPf6c6TGQh8WtLNiw
bf5d/O2w/zsjGbvDULm3dxCTr//fjg2ix3rTLRXJo5vzRWodoiHKzzM9SuUgEde3
hrNHfXlc1Xg4gNwjatoHW4LwOEzud0JFSiS/9nJXlOu8M4gJoODG7D3CWIEnjd7t
x3RfZ3uTMoKijCb11pU4cn6rsMjYSvz5l7WsfsxnUxbeSV+KnTgMxznGaZAB+mYT
ske21XLTAyWYI2eMAwsUeOtNIWcRNC9RYEIMdufJ1tru2MTNqtCNs+qEd07wWhiu
qP6cuigDnPHy2eqPKenSm12w8jK0YpNsRnv2qj+HJVP5yOp9KwbkW/1PiBusurUU
sdeyBIcNlzbExUzTsV2o1G735Gecb9hfliYkUAraAS8hrL0rfl0ylvAuDIIx8ox1
+z53XOSpDRDumKj9d+6/NC4UKMru5LbZVGgZ5mZ+/ckfS1Ea6AJvp+S+Fmb8PAUi
Xnq8jO+ZBTnYAyAaJVax4lrrcywU7Q6MMS1TAIYtBb6kmvnde+tYV+tPPhcv/Al7
2TqrBIGwtaTWZUCNKHmIdikrl6oU6RKM05TgECqMTpppLiwOorS3bMeCK5YEB6VC
ba9RaosvG1GKV8xRHvspHhiAmT8AOOTyCVks6IXJ7pXkS/fsF8wNe8s/m3UpDdqz
C773vTFxcni4RDTgEeSeYfLCSqC5CMC737jBkG2qXcVbJr5N8UzzxDvrVZhux3h1
ks0Xd5qsrzSRHPUok6KcPP9NMEQZX4J5DMwpm3bt4+rJM3jiql3UnYEVLz/dUNSb
HTw8L+QZF9toDZhzzFP0sKBHaRddDnWIHFnvV4ax+JFOYkaYMOjFYN7p6jWQBYKa
aP9YZGD3vWjQfjcvosTen5ZUpJIVyK4COFgyHLBz9TGtjnU9/KB203i9TeDLdgXp
l2zWFK50kVWHZxtNbJ/4KZNN7wKeerZzjr9MevIcgIM1D5BzrBzlG37+526GIaX1
LF3ykSkOGS0iAKMIGOhSVlSQolEp8B9EZdVK5SM19jdyqJNaSB2zibcZfEjFzDeq
dZ5ChqFfH3edlQ+uaK4oOrLOkXKJg6qQ1PUBKU1fX0Rbv/JRSO+aQxkFbM6NuarZ
5xuFFcUjOaZpcslB1W5BLQ/MO9VzCRZkuimBt3ulD2tDFWYKmyVLcUj5O7pGmEP3
Pr5QhRlR8l0Zo2T8H+q7Twxe97JEewJZfdsFoyHL8TjNROJfcKuQmVEhk4MBW3+d
trYrUM6M0Jtl0g0KVTKxAE5PKNOM17FyGEEq7Y5ry/q8sgrR5VcplmGv97Ca2NGg
h0wtQ5zfhIvtiKqUfmKHyS5FMhAuxBWP03a+gHgq24YHrMIi0MeC49Bozgy5IjK8
1/VkfvfU53SmqUUGtOf7xhCT0lqeJ0DnN2GNCAcY61tLw30M7PzxQFiWLeDX/z+/
4dzjMVJdOXu92dGo9umBM4EU0ibh6OL8r1TGhutq0XcuFAJ/F1nhrf+x8mYM3o3C
PppPUjrS5xtWXaZbuWy2C+g0HRMk8T5Q0eUH6OR6y+syzWQfksvoM+0cH4PxpbKS
2ECW2yVbDRKFcK1Egwkzy4PKPWGcimxqylUD9TpzVePC2v0vq0fpDkM49O1sibOK
WWUu/ZK4bt++cqXjUDLHbs2viWveklTYeqy+Zw67+NHzv+NoZcsmNqdh7oeJHU+G
h36h3GYKUAS1ADNu7hMF7dvkKjZAbEqclncFWVezgUCXqO2E5TcH4/TFdglDRWNl
HAYkjL+Ns5HjleWomrAvozkzAqDZAY3pvzOOSbmWcOjbrXzr1ITvixhzpcsrAd9C
E6YLfTb7OauzBKrGjWwIYWCCYRsO//egcjCog+Wl4nTAV9SIR15pdZqqaNb5Kzir
YY7fA8CaiCbvGQNSqyNrI60pRmIvUvsRYO9c1t3z75rfRf0iIT98TcTUwxMfj6Cr
EmLZBCPd9aMlEmH7JasbMsJkqG6VgTVGyfUAmlV1mj5Yjj4YpZlUTuAsX9Z1fgNy
qIrZ1iEnfZV/yzY2/jTAwlZBbRAGLYMf186CI+CezyOQTM3ThkxEIKbrdKZZaFP2
irPsW9KF4dEFMwWOh+LvBarjENa0CeYnWErKrQUAgfStZNGSsjL9nQCK5rOwxtZq
YNeMu/OknNjtpEak6rGoFHt5L8aDExMKbClmjziQNVe3tvrp1tx2ZS9UCwOxg6R+
WdklnFDDBVX3YtbBdksDQTX1HtViUICyVvGCijar8N5SiyR93zprkBF9KveqhBv+
CdrIoiPfwxb7t2vboFFMzi12LRaP5oZK0Heu6VIQel0LQ6Gs6J7EtGD4syY+E+gW
XSk6lqYYvAUyHKRmvYUENIxiv2fjKmJThrRqjFHvDsnAZQvPDCdBsJ9a9Gm80QlZ
lNYLHxkl0B8TTr+b2Qqqp1uquVGf3x3L+gkSjDLWFlj+4qQxyW6COU3usrmXv/Cv
Ouol1dYa6Kq1VuYZYjPbtztKpynuCLd9Z9SPcz60V6woMn9wf9OxeI+CsFUM4qQ8
UfH4dW5it/0z3I8l2tYc8dzLMBvqhsGnF0ffDdpXIIjInIUOVt5ykvHi1iatQeNG
y3up4Iazm0yn/6wvzj/Iuk8dDomml+e4cZkORrXq2Y9cXwAXQpzHcQ02Pjuozb+s
9IXEuwI++zbvmlvDd+uQ0LFqDxUXrdNSpRC+JiXB0YXJRtXPPJ245+m8lHCClT7g
dAicqoa4jMUg3b/YCS6/L/Iwz32ZoUD2+qaAJuuVySC5LMSzQUVd9042WmmTZPYS
0ZDNy2ZKBg9EbPdi290IO5tnu1a4uAFsj0+b1yipvJFKFF7ghPol0zaFXIlLjq6A
v73/CQXjX8wKpkNcrnRu0lyiV6aMM01f9Zes0RmW7jje6xnpaRQc3vB7WkfSI4Cp
sLWJwuAUmHd4EDAjCMQxg43aQbL621NygxqrqeDf4ZataQvupfwPxHN1HdRz/o7r
2QQCjibXSBXDjt1FlI0DyT6pUAI5FH9mz5V2R6KVl4Xn7ZoRRpVXVIztI9sPSdas
0u4mEW9AWcoTuGqnIYVW5CntTM+li8xwvvAZWMT63Q1lT+M3stqG8NhMVmc2PnXs
M0hc8aUHn2txMmBtDTUnkpLVmTaNRi2PUb4RgkeyICrTrtZ3WMBUrkdAopgyHtZC
zNcVJ8ckME8k/DPeEJyd9eluM0O1oIqpjNK050uyRZRXDAQv6DukpROPqOPa6Z4M
uxPd8rvL4yIb3NAJSZOvng14Uv8V2GceojXjy1g3DSIkNfqUqtGC77xSQ0Z2PJWk
Y+e2URxgJGqky8JmxCa58TTmsZzKoY63D12UuJaXwRfpZl18ZazvxoMMkfOU874U
1kqy3Az1cMsMLohebjS5ueubNuDFWawv1rqo4qJlb3oWHBKW3IDCSp3JMlrY69p8
t4izIXo7TXqpXlTba017r2vJAzpw24M8IkPkf+HUSuWNysBtoGe82YuIS9bWNJn0
5fxNDpaDdPrgJV70fS0ktSMujlhUPT8mMq+9+C6WSn3dnFWeLnaS8x20gD4Ra/9r
3ZIBGB4O3E11/mXWE4oyW0qIWT8IoMGeg1jnHskfu62ZGAITku32sBEEMiENkPOz
bZ8iB2kMHCuxrLGZCLmyxVUUpGP7By3sZHHdMbDlOsGhHz0RV7FrhX2FX8VKfXLJ
jPdF82OPI5/IDkjp219kPvHjLKw7n2x8SVtlDjUI/nkBorFCvTvHiHxQDT6TSfE3
eWSOKpmTtEKfcmx2/IgwlMWiLiGPKTbmh4WlLauO3Fkj+jcXeSTkJ3gqKJE2Bv6Z
mNcKjh0DpnBNVYpFPjZ5Z9xaraPuuaDGeEIjsVMdzBsl9n2vhblh2TCXd91+DZse
rw56Pg9ATcLTtexQbpmcYjbBqQ4gzMEhrsmsi2FoWSFWpiA9CTt1YEg9GSM3wYbE
mFPIY63KVnUEueG6RGHGqGvZbaimeKIDQcLBA2RKA1hFSRxoHdioS6p6vLXKPpPz
1s7UOxpyD3lVz6qBBfa7CvvmpLdZlchQUC5Yd0fSCUtCadV6pMVal8HrAMRRc2sG
pFmVlm+ioBrKE8xp5WQ3hZVsaiqt4F6SXrzNHN3uYFXfMll1WFQgDHtzR/LIxX0p
78MhbM97GhG2sT2KPW+cCc+RDGIJwioabWfex+a+Icsg/FBNo5lMzuIThHWHbJV9
SYirac08KytKj6cQa2wv0yjiR0Gbv026rmfpQvtLFe6sFX1csJFVdiqjVXtpFeQa
qJHfy57ckfTG9QBZlP/MmIWy3dFtCKboNZS84SR3x4w2cmzTSOcaQ3ql72KHsEJM
y0/7NNOhwIt3C2IT4pnW3ydVIoZQBvEMI2XvL8IschTK8xb0yEcU0/UkUgFu56DJ
pUtaUL41bCDyFp6eDnJSYhtO7y3ytWHug12acrjBvUOZOaNhS80xL0TkHmtynX1z
Mka0su/tBJdkVBYF6JJZAHvfXZ83yk9D53UzErdV7Q3QvSQtW5M6BYTrzxhnWqak
DPp3QrI68njvgaTGnEsX45PcucYYi82jWogJzGgSL7RAU4XgAmqYpaFlg5uH6JF6
LlM7S8j0fdFqzX1wj2ISc/H+f0CYWfq+nzsX2IY2bMC4dRITPHm36U9aRg7jdlAv
Kvgk+dRsuLxn+3+AkkR4r7vUdbNavKANXt6kI5BoWV9SIl/fukcSf3VGXNDc1UON
94L8IhZ0CuYa2uWdtNuuquRLADj/Bk01tCDHC8xZmHX4sh0tRRNYbpnXJbS2tymO
AKCriPUS4c9Pw1ObMkxfYRTwboUrpUy5wUWIu3PiB7kKZtYSWFgLeZsC+/vzrGQa
YhLQZy5h9h72Mnt8qHfyxUmdAi9rGZWdRL9lqW0RofRq30RABeiLUl7gDNxQudVi
61oUz3tf1PHhFa0ZZAJ/v/8YPx8GZDc5pNYhMIYMV8HFGpfTg/kpLqXKJxCG/Hbn
Z9gpLA9QLhW+ICx9BE0V51/AZeK6M68ATgyFPtrfuFr/sbhN80zAbAMgYhzdHZtW
IHcH+bFKy0bkCJnU2U2URlz7Ky5OVxG6QuHmQKdEgoXn0tEP9oJsXmMzHRcrHn+d
k3RlIY2vVCjUNQTOsVWgtlC0iaX2gU4xnPyGJSOVoRXvWxFEm5s33eS4zep/V7wR
Sa08Oa7upPMNopjRw7EfXchPDZezIL5Ll9aX+vod3n+o0iwLT+BNg5J5eazh1L1a
Eh1XwOPYM6McP6TKXtbZMruSI/0EMN465UtUtU36k3D/TzwrOsfy2Atk4dyguM93
sFwiuz79RQCGnvalXZOAVP6jQ0dCiafZEh6MpYhMKfDFUy9B6hzKzDmMMTDLUZ2S
gTCltoULXPgbCTLEtVu9eJdiOGhEMfacTKpnCcyG3TiLltQ5ssbWy3dtO363jPcA
mNtD3RGVfJCvVtWIMDhF+7gWmqUARmfOIgk2g30wVZfGU1uEXaeH3WhDvDkZYXAl
f/BIhJ7f77ZP048KuCSgHb4+w40ejRAGkHDzqjEyXe4/tYYwHrmpmj9Wk5Sp3Wok
cKdvoWMwa/MXS12QEfpStqLk8qNsMANt00VRaxAQH58grgZSURyojxBN5tH+Jl0l
BVC0NOiOR+hn69OGuZPCWaBv9Pz81V591aGAln+LNGue7izuO4afHE/xcxx+t7aE
5WZj8YFm5c913eV0fMHFxSLZqScy5C/htaZvwMpLAHC8BGGqQ+KFa6BE4enNwZ7A
6L/5f8sc4uJDMiOWithUsCjRw4Q9O1BTdbc/bbqA1Tp0+AeV7PjTu/Cz1K7CQ3ak
Q1ROQ5AYmAaLvpRrtsA1Bq4Iiimisd3PUx2IiFokY3xsjeFonOQ6LalHdCF8clyP
sdmuHlMX/P8J2aqJcmDakfDeaw9WyUeoUtJLUivh8vwpmtFsUhkoqDOKd0+uuG4v
vfTyhlntCsdCVPCYQ8Hfc8s/sMRKvmFsG6BHDvSTeDgYjuw/6SidaXeEQDG4aAPU
DQlbxmbUdNbPBTQl0wpxNrVPVoFBBbOBPcTLUwGJahnVUFkfMSvSBQxP1pZNNGHL
VjqtRIIYK1It6ZjzkspSxIVMybmbf7cAEKtFSq2Y5XCFyUKUzfBt4bShgQNLsOkg
NOZ3brB/99f4CCOtSgRWZDPKXBvtl/IbUCA/4UHltCmm40TMpU33gFgr/NeHzpvT
T+hvsRtAn4ahPMZEOU+FIZB17hmoTve2ApxYs8qRLSL1k685RM7sPnh2ti8DvneO
4do9DHSh1t5rAu8gZsBQbbv+OFhAWESJoQKwC4xDtesttQ09yba2AnRm/r2RI46K
D5R0Q653Sk4BDC6DYKbf3bsSmOQgNFia8W6J51zx4EGwho1pW54VNg/f8jFqXM8V
sPGQHfqghH9CGimDKXZ4beUTuoxld3jB25zV/3oZwd9se7d7Xbs4mIEW0DJ7sAQY
ir49VJMKkQV7wwbAZqOBVK/QqFRP84IkN+sFKISOo+PJP2LndtQbyJ0TfD8E2rB9
oSvdpumO2kM40naw3SSWk/dK6+Q9SSrJOqTWXzctRKjPzdXNL+U2Iq1hZ4Zv4DXb
FtYvQUnNLL1x01n9XZpDmIf13C5wkNX7H336Km5m9XqhznJg/qqUMkXQgi/uylQM
RkZEWY8q7i0ifx5PrxmYZ76xlI7PtyRpZV3qngG/84d6sjZWeN1lN3FGAfio8alp
eNZiYVo7yENXPJxCkxVz/dkf1G1aXda3AuC7KHsQJ1m+w2ez79EUy8O0AEB3BkyD
GfiSrbtq2Xl4WI6mnuSy+nDt6JBySLNDugrPU+tlBT9OsX+sviKCAouY8WwjhUe0
7M2B9t7Y7DobO12NA40xY/yg9AfrG2Euq4R/NMaYGi60ZQ2zsG5FC5A/9uuJOpDy
gVX9UbIOVY56PGY4vtz5eK7wgGirto4CufwhgBW7R0d5UJFwnsynOjCFPM/Vnic8
z969pwbA39HLvdTFWFEZQOuVtu80BU6PmdmM3oKw3i9FSMl/Qpxnae4qwrgQmnOf
HK1LKJG79eOmLRLmX6ucCd2Dy4D+2zvaZ3Nd2FM9afFokmz8MZeBPXm3dzdZ0Tv9
s4XvZGZ4TizfzFvzXEZBhUd1urhb+21QhSL6avtESmRxEXUyAkkL+hOLlG8VLDA5
/Aaf+qPom1KdRwY+xSi/bZj9Smn9DZyBgTzZD2QK+bXlJaJmFFBruGf/8vZJoYmT
fqNMtAMUn9LcHYSCnZu6JKD5FEAOAERpThEQT4ZKjtkUZCMheE+9GcMcnaMYKjxI
PiLkRok9z+7esVwCUsEU2gU3pTScxxSBYWiVfv7s4Sb9Ow6QLu8VSde8D+pHVxsU
eKmkho214S5JQZ+YG6SQ0XYSaB5sQU5j76ggy+sURzqANodNE7WUAYpIiYUIOIxI
zIuDy36aErbSFPJ/R2MnI3PDjlCV5r+H3GCjJY5JEjjzaPYRKIE5LnzJ/oWz//UC
3WIXLTrTt8KyBUu/4DEaKVSeJY8d9B5yORU9L5v9GL5rbMKHOvWydDGreEQcqDzm
2lawin1nN8BjVkPyrnxDAw6cltwIznAs9o3dNdYdEvOW6qmhS1ag+JqqvxobuB4z
+jTwHZOEpz4ZtGaTDTKjMPRcDSU5zbuL9VRjo008TVwYx0SJHjf4Xv/1lY2DXmDn
tqfB2SLfEYT/vY1XdKIXU3VPtKBYC81V2jZwvQwU3TMCYf7DDNODviQChJM3OZwH
F0X0i4lWvBoBjHCdWvxyK77+V1V5odMv3tklRphVNCYPCYLlGGIIS+uxCd5zH7tq
PpujzgLwS4ZkjWZ0vtNIENtvRmmRUVi6lNiY3JsKuSM0I8tOjiUaXh8InlvjiJ5K
HkjZn0X1o307Tbvwu+/rzTsHOhFUZ6AAS+sTLLWGg0UNdQankAgexyr5MZdwIFSX
8hNXCJcn0oQIoO9doIdtjJPpVjWc/Pr3o4PfwoZ44MatB/qoQ3R5JNd3nlfcvAqS
XAh7h3zyxqDeMnlY/NQ/Ys0jPzlt/s13LnBtK4JWy0RGYBmDBJxqIRkIDUuP5WTa
Mg0S6HJ/41XAwaTKs18OqdQE11PR2y/QcYY6A4ffO+iBoW0/Kw48EFd00R/MpltU
/I12XIYwvJXvAA9HNIIXh3eKs//DAih5IwWum4a3JGot1gwRIej4oZi4/r6tuZj2
AnKE9SYETIbSIvlmeNZGkB5Ei7KdlYxMyDmgyAxRJwT0nguvTGZhEIEIpnIdIWF+
bibLZlvJuxGHkclE4owfRqCmzM37Y2Sn86KPm12Iq4sgqOVv+PNLZ9OpDaW1zInT
9U45h4FvbEizVoEWMmE8rV0MwUlCrJ0WTe4kUJKTTekLyIXwV0jjCoaRC9fo6+hD
BAqsS2TAPKTdO2+1KbLVeW9hd3Vc+9Xa8Y1gy6bnpe/9j9Qb+7UTvH/X2cecGGKc
NkkHrFlKuMJYsqXn8yOyg+YWUJ+tTYqUK5FPseJ8hBq0Rr+yJ86K3jJrg10lK7Ri
vSAoV/lJq9gsqmNRQ5KIRSP9ZCA7jAlUJo6z0I43aJbPyC8twu/I1LVcE2/3AQHj
X2ypr0C7EwnxjGbSfuVaiHBmz6i514ovmnht64Z079mSZ1xmDRfBs9niFzKxACLZ
1BFsp8u/XrjSKID14GvjvbQ4E92m9BA9Ys0bTW8PQY0PkgNG6Dl5pmASwoyiZUtz
YJfnyhbnAN5mZnfWv56o9oqUvg4jg9NBtiGD2DUM0qeOghCzy1Q5ugS9+vPwOrUm
ZAoKQQyoIKGFkXjwPXMyh98cAw9iqH9VFnRglBOZ2IQ1UhY3jiV/ppL9gpaLjt18
XK0giI6j5/KWPl4ppqpqWF1dOfb7cA+vy7v46ZZkf6z3aAbjoXZ67Jesi3ilb1wy
b8AYC8GGkyoXCrRlSDv0dhxShVtwEIfB0mxI6g8qwZGjsh0x6CzwW5MxMz5ezKV4
1S14ECWPtNvVbiqdT78kEJItQKvFwEuoZKJgAOt5jtpJiJu/1sSVgDmUbqZrVy2S
HIzlG92/xzLg60ZDNYQUcawcKjfHf4S8tFDmYfUAAVnKmc0p+UwnRPaFFY3v1c6A
NbRxjxvtz55G+eCAajpK/+y/nYD//V8DI8+f/J9etR7UqMnyG5enl4GRxTH90Ku1
jI4d4zfaeNQHMpoZ6EKcdwhP+Pq2+vw9VOpIKUXRP3UdUVot677J1x7JSodw3YTW
lRcXFwADANyGXYxaE+gm5ER65YJbom/2MJr5TL9jGI+Ov2XIHHTx7ljxy24n4xz9
jD8tIktkmvuEAgtMFt+hz3V4uYdnJi0qkUs6uQftX57tb2F4kC9QXoTJ3QJ5UKKQ
7mEG57eDEZLAcW1mst4H13xSR+rLToXHaHxywR8IptgGD0x8KyJcAQy8+HhysKIE
+RsAuZRiniqMW4QDrRSHOLzDwTz2vlMS17Igv+4dCGfz6Y5gSgQhI2gJzrDOER5H
xLTtnaxFPWEWhb09uSKcmVizBvyXlIxRg2MnOKgNoFAHabFzo/OQJ85NMGabEadb
KKnFaobb1Y6Zoocqn85emqPY4f4f4suw1tio60I7r4mHZ/dE8j/mOcUNd+XSUwdr
mKFTj1U80g5X5drLRkcdu5aHNki4emAjTwmrjGsq3RsKlpIWOK5sLZLGkyocxHQX
lINg8bP+IZO0ba9qg64u+g21WpE8zFGESdOkBisIz2NVvR/dTpUUX5vgrh+8jItP
NG+G8o60m9qmgaZKMCIUIK8qx0f4A/3xh/xgg6ueW1BcBB64CMNiGOQfS9kyW4ge
wB8VgHjGj9nzVH4/aiUO54BkJDjN7nlVWJH04LQFWmJZc75aezMep3IqOhpc9n7O
zqcSH7BMD2RMoieQO0AmuzwCBjb2zUdLUD/U+UGmwKPZwPiEnR1Scx6bVh8ZbRqM
5QavS8xfA4XT/hN4AQoE4YEtG3ngn+4zdP/0a5tELlEAVT4v7A0HWGCOkn+1E8wK
qYImgD03+stPCj2vIVAxOC23I1xciQ3+jL+NZyOQS65kU1tFBosT5DfjuMkNCMD5
GyKWsekw1WxDv3N+bhB6v/vtKALFeRn8Gbb0VI2yOvKgdC81MBpadxk/tFUgpCNJ
YBUxiiflSJ9qnKrfNbKW+llIne9HC5qaDubD+o87J4bysfsHq1X0/mddxqeIvxpv
vP0mzKBwMnJ8Wm+a41FFVdH4if/8EcKO422O5Uz1ZeoogIN2YhqtGIYetH/VgukS
MIqi85xAk+ZSaE3R/LZfFdxnrv1mnsdd8w+QIP7lz/hOgG9xWA7E1un4yc+J1HVI
YIJg5zzlIyUBg+ZRrKX/hU6rlPtih6l+gOkMLlJmOj7n9osoRGVVNcU5THXOGiyO
mk25kMk3DILitcaBPAPjJmyuR69l/rrLefdATc5RFjLuorYPbgBRn0AD+XTEmDLl
hHNYoSH+SB50hr387qn/tPrJOZ4XhMC+uq48sYdCZFU9cJBFtzwL6fr9zCLCNbwe
PoNuAa3hbDfEeo5ixc0EWiILW8hV4AejqBKEWauF5y8eNZI5s+IPHf99mQTi6EaD
jZTOtIPayLGKdykZKpqvl2PqY66Qr03g/YHZkGsqVHpp/j2Vhr6shYrMqVzZRAtx
jxCuXyUNQfDi0szBIMCSwwUeoC4jBWG8Lk372h0lzlPGdKwrefpCsFgShDyKxDbF
7ddLReCHRb5xmU7T8SktQCXOB+rGpjVtjq3i2sASQikE1YLagDW5nZ3UGU575k2Z
jKYE3LvFzSrrZY/4ING/ZLry3MJ5ln3OIcPdUrPBhSKXTdvqtLBrtRF2a5hog9N4
0ktHGfiGynygBnFhth1zlPVFVZEpVSteFsBw2WlXbw4Ej79AJQGAPa+TPS1q1x/7
UFyRMnIZWqpT9Farh9bX7YoOtagNbUHkG0g8mP9Yh4O0SOJEl29cL+N+OpDpXNcA
AsLNYv3aYAfh2sW51Ux68fqoVaaQFqm1b1PvdrAKYo1NbSDHPYW7/uXHZBat1gK7
9pkTt9w1qCFrgCbFQVwJEz0fCJavl1jtyvlScp1YIgXqZMn3CFCdBS8IVj3/TsTC
H53OAZ8o3jTv/+1LjffLfUS++ZOLP0flgh0q8AqL7ONOhkulHNO/7Nw39a99xxAB
34j0DnnBDADCa4CIzrIf220jjY4AtC/Z9RT3PRnrelsUz26GhaBcQxHP932FgfkG
A+wq5dlC7GdlZJZZZJZlEpTW4JkouSgAmESFJ1GetcKQtK5ih6zOXCjRhcolp76i
BCMUiKrwikM3U8Bmn3RxAcaTYH9WXZ+roQwZ6e1xCPbU1nHVvjNmdIZfH2S+8VHl
7Jkc1rQm0bGG9JHLr8Xl040GXFaIs9EZR3Xk9Nyp5Sr3b+dZQU6+L6RLoltYSrSe
mAcQK11OgaM7vyUCoAmO0RxnEJJmxpcE8Z/ngv8MkEboZx/qjT5xryWdjTkZtJEO
T0oipQzqfwxXpqiuuEoAQROWSL+8Es3GsIUAan/8ObOeLPF9hEGMa9mfdcw5a8F9
4EXKgeKInISf0J6xamBe0tBygJpI+0jqeu6IYKMKlTTG4vY8ktf17WvVrln0KeQ/
GYOHMl0tJ88KHAL7PXY6RJX+JMk2vEtZbaJsquQ5QK4kNB+7yZapKea6kXbm9xw9
RtoBLHXy6Kzw7XClcibsfmwO+YbJgJfGpnB/eLXQoFxTMYnIYdkjqFOeD2Y6WRQG
v0q3BXNKJ4uyMSAKIQHPFPI825DgEE0EcsE9uwP4La/M3tedtIIY3FWgEX280FUy
dozdYtFfTEUoltiGFRWhijVbOtFyOwnYJnHWHSzcu3qaxvIak7I7inVzsZwhcsKv
NEXUaeaMIKLVsKgL6fzKUSqCyqjeaWmtLLqydTr3oSNQANHvbL7fwbG0dm5V2gi+
+4NbXD38MYmIGaaF9ag71+NGhdymJZZAs5vrwEZXHHu3tftGha+kNWu1Yvd7qLGp
pszPRjrCV7W2N8xrtZX9A1HTmSTv93YsEPTKyNeeRZv0cB+APZqQlLXwhsOaiN1M
tueWYjrD657ENmu2QgwbQRjUZwFVA88nxmkBapy8Z56y2lztqk+zW3/YqbUmJBLH
wqbPMEcrjihG8zh5n3kf7gR3qNQblWFNBsjVzuV2ubj1OrfgTIe/NtkcySqq8XTM
KKkE1zinlbUNt2VL/zBv3WTf6ZEUVTVChzhbChd+9VozBMA1MYJ4c30ShoBx+xRx
lfy2gt5yJ/NMtCEIThi1YFr2GLquGIlSDeGRTH0BgGPbkTz2rNmq0ggKhttrS6F5
Leyif/69BhERVIbt6ufgZ1fHHH8OsCe592arC7plVu6AV1nQ/rGjqPp+PtR8L+7z
ZFORdTLsY20+xh83FHB+MOCvoKQnqIX+HxgUDq9ZghnGUxW2OBmZY7Nbxg6+Ro/3
TkEqayxAEPZl0Z9IpDxU+CssMjXw5RMojpJR+XIUCFfMiqTqxaR0PjvPt9kwS9pj
OitjsOT1BnRVff4lQYujI35F/3VuqZEURw/yRDfJcg0/8NDF39KAkA54fI2ATPGC
eB1WHtdznEOoASoD+mItpQVMNjWnXDyK19L4j6pYVwRslnjDXgK+vw4sHUHqh48z
7BkCCI52qy0isTrtPW0JDU6b/MQaPrE8eT/C5SXEOPUTUTmYIE1tvQ5v8F1QM5ox
MZgT1ALJ8IKpjy25lrFUyzPBgk3UEFQxVMdxJFjgCWCEsQtlQb3qIt1RXCUosaRP
8Er4QqbqziqPiEYUZWInoJRsXhObEcTt2hSUHV/wW/vtEZnJddg5IB2dIJXibaLV
1FhjJhwhxX9rNcS/nH9x46FCyKcHNPVCrKTQvcwU8HdcZctiuehzYmiXEmeSej/l
vJCtLqnF8g5CO/n2F+EixSzIzvyzCRapwwfsyRCtEkFM8tHa+BqFSUZqOm/e1jjf
gW1wAWMnbKbWqkpLM1DJnoQoKAiCYvbxODXOepzOLMCBy8s3EkTkRLRyrQIx0aH1
kh0k7LoCEXzNvSadKhsTG9CbWPdhCCPO/P70XflCHJ47qQvPnwfngf3PpcyoBaT6
qvM8Xo74movNByrWsDI7Vq/65WnDeWD2oCDp14kwlre7Hmac63jDwZJoKpdyuNje
Z8G4rXS8K18IXVfE1AlQ77dYPdrCH84IOyjj67kTwuTzO55zeEWdYanvPyMsnYjl
yYVSyUZR5lzPkNfTSyPH+UvwYmVfz7bx5xt0INW4qSym153Xh4IfKgfXTOqAFrfA
pl9K60JeyyR7CHm0TnFVc+Zz7SVPzA7IoCGF9RlBcRzYic8w+QzIs9rH2KG1nNy+
sHvXMp+LUE+XU9G/J221M0U7cMh/YsEjbLbOfBDikv1KE4trHSkZngEvLEuhlSIm
s2N46HyNwWu22mI7JEy7wibc//9ZT2KB7cqfEz0ukQ9Bw0rFlyOa6BnZrYNUVhSn
y5uPEUzx9eAh8LcF4z1+xjurkbyoHWMQpVqk+HzPIU1PDiALY/PUlFzxXOcYOdkp
QB/3uXWm70qCDYO1zt5xmVwSniAfgVTXviMbDfU/R465zoj2rSSonpTLLJQlfiUa
MORBMsAHl3tKY/RW+iefm+VgJDiphFythPa7M/6IbfQ+yCEUoDiCJ+7TspqJoNWa
r/fZuu6PDuYUYVbcIpS/STavzy7a+rY+K/f4UZlmo7NH0a8ySGeYQ9YWnAxKvqhw
tvnbdo2crRTuJAmzBG5Go1iNUgE82hc98s6TjI6KLosBe5IxetVVM4Kzvy7t/dVi
n+UUpft9UgGZYpd5Rrf5JogUX0pu72m9s6j2thNskBv6OIefJi3fgCle5dxabIVp
ptUPwGmGef25WZfbAY8EIg/7hEU1mho5QKDUR+n1kPGsKknq/hPNGA+ZPVwCWEgw
xvwQgtz+UdlAzPvByqnm6tqWckfuSvNiyV6ZyYUrgPbVmDb8ho6SIoM4yutbQPyy
VQiB5uDuP1yt8mOIReo8xgeJZURs22Gn24KhZ1inIodywDjzsaZYPVB1EIGDeKPo
dWNdSBAlEv90Wsx+bQDj2jBqVC5XSaCzYykdhKO+531QEO7t1/KEIPMnpVZaN5II
mzIqjSBqrYGO5WYLQ/x5cFcZlnJBnVGvOsMKNxpTYM3gMLs43jp6jvj/DK5eqgQy
nat8IbUdCGDW2EsF9OEt5ty1+qbXsxMEuw061phWgoxcg1d3jnFZPnz+CVYmfzZb
MNO+d5fUdN48f81yrnj3M1qlJVLVEcQd2YGcxiwBhbCtPSQ2cg1HSkumcf34Y6+g
6Qrvrbg/lfaKb8ZI+n0KtAXO1UxlLwcyrYNIapm6URbgIUTk/7UxBcqs+bvhRrHi
KuWU1Yk93CdCmIli523IX0tg/yVn72SFXXRYF5YJvspS9XE0qfjX3KN+UFTjRHeT
yGzc321Pr3Ulxie2gh0ZVZhHPzcJPDPTmr0/i3MI+4koVYG4wZ3pS7c/gZZJPKvP
Jjkptr5Jfd02lAwdyI3amrl4ORn5LkMOkbbWrY+dM/nFf0xHp8vPHjhi6kqeIgDn
qHCajvRZREuvgk/inNp6EtlNuItX3k27Q9ubD/QT+Z5QGTH436KiDOEBvwOswNO3
rvVT6vq6ANGZHhC0/hJm+gAYDki9EIYjh2mVAQ7Ahzwfiyu1Zw7NvaSoGO/cjXjh
ImX0a55nwjHcPbc/esD8FspgXR4OJ3rBTN56rKrAZOJhJPkPwNljRSy7PDgkYv4i
Hi6dBUrvvT/lAO6DxVAIzDvP9qDcm0ERILXKSGHIPIkX2X7ocXcNRyuu+Vrf27bc
VRJyMdHCCtD9L9hcuGecosNPsc+yvVXOC6GSTl0p4QBvaKlGhjnIUaP8BOqNPTHJ
ltCnuzYCd1UKLh3+LFhBd7kcSRwmEcuQSPQzRlKzL/upPEqtxnFintBahG//i1w2
48LKv9q6dzVgriTT5+S0y82++DItEs9ETiShwuRFRJt9thscAPf13SN+CDpgbMhe
agKD8/pflFnZKsdUsl/7SWWXThDP9gVNj1A+HF0kke1NomzEuI7g0UxDDxrO9gR1
4r+s30TcDY+whLEAP6tAWdxv6vWqD6eoKYra4x+So0EoRLb7/bw4yMAPfv3kNht1
Lxkji+K05E2TVx/gLOCHz6PZpr1ezBWQ1LiCNniENjEFP0QEWYqMv+RlRt6AAawB
F2aEWqKmVwYkS4C0bFCDKSesDPONb1wa+KzmMLuJEKd6trtO4WSG58yt5a8uozqg
Lx5RnHI+rVdLPT/ko+kjdjHrJLF17csZN2ggGJ0tt7bzuHbteBZBGG5bRDkJSjGN
3R8MS43t8I4GB8FctbBQZyryb8RqNBOnuf+VyPoigzBPx8iYIwxeWWe8hn5H1Pgk
g2gwWA2lKdmXiTtASEanHDeOgMwxncZW+PML4oUY79D4ZllYYgGmb9OOQcHTEczO
7hXrr7pJ7f7c7WyNwcr5GgV8yPvOrs5HblyImym/g8xC/CzYJvmNaHkYnrH7/895
bptdd76OkFddoBAebW1AFm/wBLSKJfs7kQPy8ToyJ2ckB/GdBxJnATLdOr+rzo7U
HkPnaEGKK+Xp8KOGdH77eHlPO8id7VGeZ/lfFvn3jHs5wfQFqi6UFxxbUSj4xLXH
PLKw512NOG0gYXgAOAjQP0K0pkkQfO/G5mp3Q8SmOXugSZ5OjAe1BX5s2HiIvFQW
Q7q8wdflVT66YyLqFfQw0isIGrk1bDVlYmwtSu6iClHHFcIfkbsGWnqFID5pjas3
WDGZiUl8KMFJfMpoxvIqdLSoKjDOhjFWKPOLy/6qnt9jZQzsqA/SvVKfPsp7tm+E
at3lRgLTVAWL/l16o64yLe7zb3it5hE7dRjLMzTvnARNIEflZPvSoSOptecGY+tF
vJBUYTB9iB4x+Dl9V/JL8kUX4VrZs8bQRovpxtiPOYTfaQ6GSh84XVm3fWN1TDrT
9q55h0XziZJf7EXDgsO4eXAcrVe/nWUIY0oqym9iN8O8nQs+E/GnDSQAdkY3Cotk
pOCNmDkHZ1mw/Db2Dqu8D1ZE8xZrpwM9XAcTm6ImJBUbM4AWRCLasIKFgq9Tv78C
bXrzOBj0352DKQOXQluW5YaLkNPKo+5yZMVW70yhOl5EPJieK2g6CJQgSdB+Yjcl
Zt4OxkqE7B1cGVuGC/H7x7Ed44OTU1g8ci/rO9rV8R9xb/tiuvDKmHOacJIhdlxY
xTXuFWt/BSvjCJe55Asbgnh+HgaUbc6tUYE6Ibk/ohzsAtL3ZQEtr9gCIQJ17Q+Z
jbETwLVWjsvcwoSt6ZjHhegE30rBf8yDX/Bd+az8IX1jmUWO3SoDdP+zRf8TSMir
gtgOSQfJiWvuKXuXjbuexcNvR7Nl0aqZOleG0LzFQfvMCiUvpRHhOUN6E4O7lso6
vbWI2JhfPpEbLPN8oBv3uyH9UogMTrehkxovQyA1qh6HxiaP/uVuMFABUaGEAMNn
sO4o4vd2pm5WJOZZ+f7Yvoj9xH0Ci6zxv4z0dc5ybXciFvstujaRoSEWIpTfxK20
OBhS7/3FxylUHWwf/L+lTcMyo9vkDLumIwK1TXVnpGtjnEl1bqtd5SvAdzFwD9ns
znda92zmSpSlQtu16GYWMVoaly0POkLF4x3lNHg5l8GWFFnLTNlZO48gtyXYSs0f
IgdowfFxN40UBWHpTSjMwvY4AqX3remSxIstFLJrXeI4DAtvMPheCCL2C7BDZQ+M
PpcI4kLHDCQgzR35hnKJwKGhiQMmb4JBeehywikkgvkk0TjZ9jKxne3XE7coDI6q
PD2SWYZM6s8XG4/b+OPOoICFycc8DTrQYXCOXEVyiIdEdqjZyI2ooe8UgYCXfpYK
aSnbO3sOJ1A+znm1rGgA+JqtObYl6nFQFB5KM1jYJ+MR9zc1+l7YB8Dw5hhFS0HX
VZ21hM8VcpbQyen866lj9Oux/WcOyDJfLjgJvrqkKrhGSYx/p18BKbZWOw4yLomy
akOFX3H8OFAv7BAXGkt6AKj0d+FZttvgneSTpu49mC4bEoVmD6cCOTi6UhFb+s0n
H5FOhgOQzNeVX9aM/JUeIsiopxsuerAf/ID85yEIkVZulgLMUoM+8hIeuhIEVmsi
WDL5bX1kVysxBuoxPhHQtG8AlcnausoVCEkMWJ9ifPV7MglXpEtPOsovSRrns0RR
EUk3Qi8txqAYxPMTruk0tCZj12X+OmBZ0V2NrEQTqzmYVPKqKpQqUc4FHubPntjZ
5RNYKE+j1XZ0B7xHUe7cTNzfPACwdT53M+Sm7pTVqP0Obc4X9ChqLAqRqWmpqDN1
tb9FYtXwx2D5HVGgXFtSiDX9cR1fsVvXTUgGxF1y+FAafAgMQuWBSfgWj64dbU1U
C91PFi5/OFfp9Rg0s7JmAgc+K3g9p/uM3SxD/myfmGvrdkxUnyz7c7pzDVqPVDhe
LGfIKSJrnJalnbtd4gu7mglSm1Ujy7iOwc2gyzmSlfHO3tqElzLC4C2DeAF+Ml2M
z3J3g7ytlolwxaUhnxAHokCNUDzFmTIxb/4WYzm4cNlHSC8b6loEs9ZR06jVAoYY
28m+9dTxB6i2DV1Q8DMC8Cs+gM3q1XfG3xPR46n5ZREwUTR0kY/xL3ylBoTodmir
PPDUmSUnA9nRhxFZVHm3WHAKi0UC+oGDtlRZtna9eZMytvd/MCjonc+irHd7ICWI
a0u2niZUxbLa1Acy7WrgUXLZiwTZCsgNl+uqBerTvrmBuffopJLV+Gbk4Ju2Tm8b
d1NtdtflIp8Qk5G09f4uQrD5soKqoLHhU1/ZtNUtIbebqs9movFSg0XnoXL856vO
P2sh4H6Ka+1scwyYgIjhdPEwVSQ4PPTWsF4xsmmtkQy45GTPvYJKiH2yHb+qaaDY
tG3H9brNgOG9mmRopNDXw2HzuGio+SS1uEVueFHqmBi8LPPXsMRhhGZsshjv+otd
jO0PswH3xC3jMmodPnjFTfxTgpovZbpyNmOFLEk5EPC+mWOyWv2rElbryLFjPFg5
OsdldW2qlmGgPquZgVrfBwGO+ZCo1Msm45cgoMYj8Q7Cow2J55pxOmGWCtUY3Wmk
nQsEphUSk1HvmWURPzj9KCVqSKRnprwroPo48x0KIJN/EHGSq/t5Kpgx6LRgnsp9
Lsl5wt5DEb2i9OuztIA64SeReLht9XtCF9VKIeH0WX8kHsX4YZTsB+kgbtFVp3wh
25wiiCk6yA6DGI6noL3HrqaXo3hYS94zFMO/s6TqQ/yXu3BDR0eIEiTfeWDKwNnB
SEeCamXseQGtWQ+d9K+YWqsbooy4NMEt22b+DaVKXejA5bvNQFNZdch28H1NTDaB
EddnwhSNhaiNssA3Iin0EKQrmb+5XwcsKOI5rkwuW8qAge61/NtRuc/gnYIF65TV
mO+qhRc7/pWAfF7Dcc4xZL/bEATM3MiHXnRouNO/cQaF6OkV0nnGpxC16DB0jRas
ULvKP7FgEMoR7aSaGCzEeuQ5lAissq6BOGHkzNFE9aoQf3F67KtoEOZPz4hmaLY7
zSQY/nDui9eW8wgJ2ZMx9d6Xk82NdqNDjdjQLwQ/keuvlWc1J/DRL0uhOrfuW5BJ
6tgc+1gpWTiNqifzcxq+EI9MAa5WyJwDrVxzQdK/K89EMdRnj/eKeQD+/ecmV7x5
lpDMtPDU79iIWMdfGYbn2cErJlbDNTMuC52F6UfD7zE01yBjCAGIalXLWCCe9GWF
O9ScvQPdGyx5pLAmpLQ1qkPm0BfioTG45RQIItfq2jnXwS+knkrNPMN/v+dnaWby
g2RgaLX9Zzgsttw6GAAczlh0DiIEHdH315QKeSn82WAu8xtXL+3tp2B+YAiEwZiv
d/3WlJyZ919GV40BVUzTCKDglvVNttvguWo/Xs69sBE8l2RJMxlVU7dyC56Iz7B9
lqMrQT31xDCGM0i0tTMYKYE7o5ZyDVVQa9fPVquqrK3pIqqN4SGZM7BBq2sKwv63
feOqHi6Gxj08/TOzoPpIpDLlGIyd2M2iVkTS5A8ZCHf/pIwJbixN+Ir4Pyzh0EEi
evdhYL+cbqxjZ1zWpPkEwnfUkwt9ZLTrWObM591qS9SsL+JqzGjRxVVUR8/3upAt
uAfT9LSSPI53dIwXDNubdEqETiN/p1/hnI6oo7SpsXwUF1pYKdEZvvQcu8WH45BP
B0AV8YzDKnc7vdpnbpXqOvqZZXiSHMR17bwUa6oBuhAG2KScrGh1knR7ose8i//M
f2ex2Vjgp0mlirGMjNZ2kWH80OFWPXxs3Ljw8dqSCWWQILnbMziVaa1d33G0PxZ1
Og1eW6MAx5v8/WIVIJCULZloAiD80azWqiOH8M+wKNeXfNngxZpfJWFfJA4Ktcyk
o9lLvDGTs7u4rjsiQl3nb0zwTET8W1j5Dk9IXOePE+eXu+d+fu4U65uB73CGKCUs
Ptsy9H9xgm7zg2BifrrvBGCbvaKTy7JC9Nix3RZmAu+i7Lkqo8WUM+/XMxsIH67l
IZlEKM4kK8J/8+A3PJ+XR4rv/8AhyhNy5ThkxID4a6sK0/LNiE19J3DM+1CYD0Vb
o7L4O0IJsRZqJ7vg9gdvVC13E3LIv/Bv46okWJ1iyzHhjI6S72GQ1CvnItmzb+lk
Zw1jpSw6/7DI7VcF+TxPbRmWBo3vKhwtKh/6opqPE7mjbB5dPQOBlgaDjBVmF/ft
5Ku1Jbj36GQ9sEJ0UjdnpwZgzO8AObofa+9tfbAKqAgWsyJhxtk04GP8VY5C2Kp4
qJmW+/dGu6YjYpeaFtfxPt0B0dBF3HKP8uo/0W3wUIClFBPUZXqQiI4eme1/gTuD
Y3QLZzn09uBnvUg8CkvAnlest9iOyHT+/KW3C5HDLxfYpZtHzj4IehUwuKaDBRQO
Iycb+deryY/XmRYlPOm8vsTT5V+uIs44IoQpqkNsMPQGPuCSdPZoCs/Hoh3wWPTo
8xOuKXm8tEzQ/0YLoEZWHcmk8qCp5tSeKT1tCLFaWIjsbpucl2TMjcr9FoajYlFA
0I/KLz+9Ayj/1nxG73+Irs5dKTl5tB8yyvSCb3Wsjto+NmGyoqLka0DvZZpvjzmI
7G7m8LXrNb+q4yYrMr76KKmQdgzVJQLXW7URKvLZSYOPQscmMfAlRWpX6iM83JzY
1DJElD4gBGrqzsHKnU35qtZ/FU5/N2pUZANYr1FPY+fag9i00lcdOlQS7Lk+prnH
s4yuGSy6FgXFNZBzeP7sYAjSXZgDApADzbCSLrh1N2Nt6xtP9XgqzoeExeyb++/o
fUL4esD0olxgkh826iuBOC/diLcPmQVf1nM6acWMGcbhXsKpHzXNdegMcDfWOfDC
9Je0XHj5XWxpOjXePd+/pwyG5dY4OHk1wC5uBAzdr7budAzobRKJ/r5w8ZW/PJRZ
698rfr4Xgxe520XQnbcXKblcHZ2CORS1KwOdoV80P1GK2H/2mefWzK3F04OOLXHf
aMIAw1bJsAc1mOy2FgT/WebRnB0ARh8A4mfHkznYuEIW0CJRSjJDZofZdnGlOoUH
o6a8CwvunrnLkSr98MP7m48dJBjO7JXsGACx6bWcPIieI2gEa9xnbi5PQSZb5ubC
uh+zuRuKD+yHuGCxTQpvSC/u3qrC3iZRt3nNmiFDQeX8zJVqkV+zhwQOKFfjkGlb
O7/XwAS0GWuv9PD0i+YYefCA3rTJpKfNLUpUH9AjVHrC60Ugs1WLn56QLjumUXRX
/HYKGv/Ux0rOCyXccY2oKnAST2k8YC6fqoH6tDKPZl/BaBMjyTKTxZUSQA7VVQr5
PaouG8gKWmConQK8cOpMgW+e632iVpZ/Y/VLaoIT1xzjKUBQEvUGa8CLDk/ijKO6
GPnPqvgILETVy7bNws3LBwNUMnZOtQg8i1Yr6b2IMY/2pJ4py8GanP5d4SJh7I5l
qKUCqPnflSUFi70wl4JxWpjVy+JNHXgQVLdThX0tEbmP+fvgKGVDk9apM53NBU56
1ToyEiIqbkacylACS46mGkEPCY3P8smKWQ9609spCk5wG+76rbX+7B+zNaPl0RO8
K0o7+DnxF3qPcesS4D3xuhVXdFH8CFdZs7/uA3A+EzvMaJ9yTjdOqOzSD6aZDDG4
DunotpPen6TNjbK/81vUpWSDsOsaeO2fquDJynECh1gLq9FcKq8fZ7BaF4bo6T2/
drKDznSoQ6XMopqZ73gt3YOUNQaA7yUbfNEBQjtToPwB3+OiYV1nNaEXV+C/wi0J
3m+n6Dd6uKxTuNKymjVfM92AHb3qEOtIB+Ri6x6nZhq/6aWaJ8QdoSH0zwjNOyJE
BfqUl/771zTiITkwsH4bZZdLYyAD/IBAusrVrDQl3HVvEHY0bvbBF/S4e/s+oLSb
cU6o3x/1sega42CQYZwvaJu6opz3JfQdhqaW4Mc9GxlETNKoc5n8pz7f8OKgFhWf
YEwPYm1nP/EY4AB05eNLKnz6XYyUOdgLe+nLbcjq8eV6AGKzHVtqMe6VBYUKvNGv
68cbYxmEeVd7io0UqX8M/yzjnOVpVgcrbCUX//yMImUCLMQlIK0PF0GG7Qpo94Yn
xa+0/oxmYHGY25Cn95IESqgsDP9Qck+iQs0JlYl871mOjhqRuIcCB5HUjF2w14wI
FfotxvVkOPaahtzgK0/WnbCvoVggGzPEEs1Czal/S8CIZZZhiX6MrEk71/SKY2Rt
KialaYg3OigoELt7kv2QTsCBIbJZGuZ90U+nvWyK7SICcQhYagmvLa+g/KKITsh7
4S6SlFGyNpYJlU3Dbb9RF/cihZ0XXPVQzwveMAS7oaa6mwu5jMbVykUR7OXlBmcy
xd1rAyDBIZdnUTkpLI305OJ6v/0Tug7Y3Xsel3iusNnS20mtNmsPeeNRw7GpPRh/
miAGm9HxUdjmvbOPPdudqYwoRDznQQjTj2XaUEUm/dpMCdd9M4QotV3p+P+72OH2
dKaA99hw6LWeou0CX8yG2tz42Md7TMyXddbCproolbSRZWBiadXrcV5+FQK8UjXN
vmtti/cmqKIjAULBH54I3K9VAehPOmJLsCDeFH7dDpIE3aFRVvthJ9Bnlkav/XNk
RTOOr+MFZ9swaoKPNpwIZXcpLPWSSOQYVZiUcUmV3upUQsUkI4Nwx7Rragz7kPeN
mik7s4BZJCaL8qrRYWeUidMnup80ndmyMTnlPL5OZ4uzVGJZvnFzDfWb6xMUx4om
jXEFoKzz89pNi0I0cUADHf6tf8UahwU89cR4ulx5xkkA2wM4M92YvQ1e8yC8sF2P
MRCftm5S4MpXoLTftvPArV/9LGXJ1VI4DmpKYCA8N/fvRBoqXegXElS4XwNTbDOW
Yea1hpC8orV2etSo6r4jqeFm94rTDN1s2yFWW/pDemN3AlSRa3E0xlVgTIzNMjXq
hJXiPjSdAwsczQQq2lWChb97/irrV8NCi5lhrmay7ECD7ji8AiCfuFLfAQeUniYk
EjOZg30kAfXPPIa1uqOEb/5qVMZ9ihjqN6ZaT8qg3Fvag+p7MIWfzozAJTDNXa0T
pYxwhAZpVr93/VAVJcuOTneMg8H241NWm8V/2pdWgpSEtRNpiaVSaRRpmYvtU/ED
jkYdh2iltjJwk6UvBeVXZTLsf/l8JObHVRS8is5iJGleyyNzSiTuo6M5J9yQm089
NZqXFhpme+cbYSE/ijARnHLq2whVkYiHoB//1Agc72DQ9sukH1FbQhUEJED1ya3D
5CJhd6KI7l5kuvTbprWgdZ1gnzjs5bT/mUD1+puETxT8sh3S1H1ZF98H8Rt+v76o
DW2kIboXmFJpJHXSD9buSMJEY4nj+maSuNh8tdWZ1h2ia8b7xZANRdFdaLwdsqGK
F7pGuuYz/sl5Uz2yXwcVIdPriw/lPhfRNlgbZnHTsDha+846kxfNwMVGNRfxC3Hu
0I8/i1bGwZfYJgG4Es8WjkLICN53tvdVmJisjP4DjBNVAu4zckHaJFletMifLvnF
InrbV5jA/3GQX1nWxylYuIQZtd8IRsqPN8T+aPMtwmndyuanzzsD25bI5hAldMQm
DWhnfqHJRGcWthiqQRe7KEUhqBKD8HizPgfnhMrs8V4Apmjx47wkCcjMmlaejy/a
29xs+CBr7glhQji8WYphfJ8AWN3Amruvj9KbqWPZXineg6u9V46gXFudzVKogLG9
iNAw1+QjojOuD+6y18tMRL/o/f1MWVSLEVNycbGuXI6tsXaX5QxiTASV54sLLORL
NS0ISpQkFhGkkNJzEKvENGxeoY0zPvfuPc17N+Bo3WNvnDo78VkLjX67KSFoZY50
haPeefeRecdjI0p2nx37qHO59OBxZapa17anQJ4EJhPT7R+OAoaxmOV9Jn44ni+Q
UTReCKEBxAPgnCueJ+h+jfGSbbYJzDBVYh4uu5XA5QD/anUJKIttSxyruFMK2gTC
djHp4IlMviuA5Xr/Ptyh1UCMamoIs3roi1eIN1KIyyHLOg95qeofcTlx0Sqw6xzJ
WaBX54gncF2WfcTZ0e240U4IUxjCjRHCUgRu6Fb1u2mj6jk4OS0E3YgPRaLdhCZb
AK4dAPITpAZYZL0BxWL7fKoIha75i0OGqris85ODr1r8Xul/PKlDmXZ2Cd+KQ05+
B8oG9Ynt8zvm/kHOJ+IBn9PZ122uf+pNXj1ze3v7Wziu43rGxj/PdqJUL8ED+RCY
qp/oLlG2srSJ6YuV0gWnPyf37U8EPE1teGvOhWXInfoEI503CPaQS0GdKfK54O3y
z3IE0VqS3bwJiYqWQspi5eFNU0geSvRZTbAu5VbDFsxpGjuz0T89gXNidmcDqDff
yz7tU3llWFokiiwKXAEl7gv0bGH5Qhz/n6fEo+k5zHMcLwJqJbC+04eEw38OBOHe
gNouFcGuePlO0CClPrLvnK44Zl9IA2YDcWZk72lLKtKR75nZrlYn/K37215Brsp1
FnXnL7FaLXrm1qr6YtbUrwtNm31OftqtMSy47QnwP2mluVCkbFpKe3WJ056RkMYT
1bsYO0D6f04q8owjorB8wyKV4fPLfU5Qi3cBbL72EGV1oyGx6WxniaTux4zbMfos
zlxMZqVLzurzkhwcyAtmmg8BtBwai8lU877B+mxGgpqOQJ6lTnRb3cZFRrPTRUoG
hatyDo5oww/7d28wWxdvIzPyIqgGt8faWfi3vDc1/OW1dV/0MtDbv401GEHBzqg9
bgdpcaSYLf1jsJFZQN5cvj3s7AaBjxE8DqAZ4Gz95NZuDNjxNuZagqH9PKoWYpfs
hvUgK8lFJw0wmFEz8aeFC9LEFyBLnBL+JSUkSzf1jp/IAtuxuuiVxSrUFX97ItIT
GMCTkGuQHRDycdu+6C6UWpTYhwSjG33aGUeZhZ8F+8r4Mdzz28Oebvk0I/oWK9IZ
VRUdJZ/0fucXo2/QL04ydVti7XBX81bsMMQWYLrMmyREbSlzNTFI7uiKSMDdUL1y
8y6256gy7IPhsnA+ZWwa2dSpuPTVtY5PZczMTl+X/7Ol+l+wiE6ngPvMRsYYdF5k
4l37/+Vk+uG9ccIcwQx442mj9AZwp3n7APBTz0OtJeznd0r0QurmOog+zhm3dVks
TaG3Rer0MnGxQtiTg6ixHPFUTu3q1V3U/7A1fExjuGhdwmxLEv/K/h0G+C/JFODk
KD/YKP0m3nZmjMe1Zee7FJrTmvOZ7l8K8beEGPsF+u5ld+WC64Gt4S9g1LR+Gb1y
Gk7NRj6+aeROlxV1uzaDNTfp/kD836ZPE6bcKPhK2t3bR5oCwVGbWnQmhVLhShwr
qWiYN6Go554ACy52oOmD6P6Ft/EcPARlyG3btU5F+fMcA0Rm2HUgBIujkoEuxpHc
K9EmhrFsqLH+k9kCbi2LWiZ+dB0rnuuy0Nx0ZgwUyZ6qB/2KXOKxr3Tw2YUyP7L4
8GrCk8ckMpdtjM9EFQASyrjNU0og5dn119CAKgjMgeQnw39R5Q0zZw3Axrjl59Mh
eU+AL8GzcZF6/NbhTImnSjsQUdF3Zi8Pem0fq/H5n+AwYH/fXikf83x0ERwkvxKU
wO16p2Gn7/m9FEo02XSLjpfUEZtXMofFi24U2g5CUkYYh5clpYegjLdQhnQkFtzM
bGm7ACqtTbsztRd5grjfvlUI7NKtUoYnncvCuybtL92tCPDz/SS2EMUotlexIkbs
wjnp2AiHq/h+x0PCW+9v694Yo99JmoJy8qmhVfCOhBy1/sVRYq0As7p5QPII8wjC
jEPBw9PuIOHApCsQkYxOWU8cy1m5QMbhybRzBRu74EOAy39XbJGWCvDNYdgnCjcl
GQP2T7iRM8UIaiQG8/4esxluTti8CJNUMFHZ27/6yddIHbIx73/o4i/2QYLfi8Kk
BIwWVHb1kxlNyyBjvq4gLG7MwBVtcwErSGUthOr5I1hQGwk6uVhh2niPu1tNcR/L
HklK54cEwnaW8Ltb7mXcsdU7pspDd8heolLgD0u5W7xkrVxL5bcN8xjbYdf5cmS8
Al5T57fPadpzVHgS1uArTjii7nVuUtqDitU6FMjErsI8fsblZoB1v5GcOP0olk7d
bCOFBszbg6Qw3k3mCq+UIyLMnSDR2A9pB0KO+Cin9IQ5ohZI18GKjcUNzycJnCGz
kvJrt4q2jrLWt74bn3+S6RSUfmKOoMhW31SMICuMHWv3PDcT+u5KtfJEce1tsLyk
ECiNQSj3TJMjQrMu0Dv+KpMyyYR/sbQVjOMg/ZFEQekqaVtRqrEhtRRvWq2tMiTL
BZOwOYARLXvfbjoM/BXwF0M4lZzFbYBZQPGERfEZpSSV1hArsGcXgLjSshKEzxOr
b+1z15MiC0/8UpkePW02eU+Q8TvJg3ssZ1woYYwE1wNanSp8RW+I49T2cIucP1q8
U/Vlf/TXz1H/w3vEe52jhZrZJypaxY1uuFlRXcBZeekB+QWXszcKVZRgFCw7HSdr
UtIaYAHx0ON8gB+jx11A8Rn3FzMgF8u3ajcyQJWbH9sacIhMdUgkrt0ksHHyAnz9
B/A7x0y3K3L6SNu+DvTfOzJxRY2ieJEkutoKuswMfzmAukTwAa6AcmqN445mKH5N
Zu3L9B30LoSM4461uN9QMiiA/9bCu49UO4/fXvBVO9m7DoOLzJGH6gg5ex3NGsVt
Ny7jdG95rJ7GEytvmJRnjzukKKFXe5IPNZFGhYA72CZ8ujZclF4BLMt2cvrLb7ar
fdDhgtHCkVoKXJqCXeRgxvdCM4cwP79RlH+lnlF+G0SJViiWNEAuTw/tgY9aJ4SE
DurX4jomorJNOR5UmBNlfTmYbc7os7C1fDJzoeEqX/jUZLiqWg91eqMXroKAHpnx
JQrAFualA98TKZSnWP4qNoEHZWMXa/xFJQEIwgOX30OOpHFUXwiOnSWCTcRwpmj6
9e/18asBDXB/oEBypLcSFnVZabdS2cAYR+qvYMeOa3tzlbzrThK5RT3J03BBG9uA
dyKDS53w7Bqjx+h+jmwbYhYLtrbKTxhpP9CCisqEOoHXxubyxd5m/Kz1k5OdR9GE
hPVVWyGCHQrZGzPxY+NvKswNEayTXwSu7r6LAgxfmbQeN0uGfLjTq2srubaye6Up
ReW6reGYwzJ0eqZnE188bbMKb1nRLhMOmB8Ti6jXTJxENKWKycpzAlDD6LXeP8zR
hM1TO72hTAtvHBGips6fIZKh6cbOmxnG88p+Fu2UtiOm4Q4Jq8XEezO4Sco+UGUR
DqAgSGAu51Ee/cJpXR+uN5vWojWNlnJLp6xImi/9lEIgtAtoJuemZOmviiQt5ONZ
Ocs4+fPukz+lfJFLXCcbplgva728TnUoetmYG9c0MEOuzmPk+yXGaQFDHybdJfk6
EXVIHgXaXgZmtt58OpTvTCsayk62ld52LHpYi/GMvjy9zhjDeYyvAWg2p8tsM6Hz
bPXtJDHYKiYCeJojjgmmJBbCSYvX/bAYT+4BDfq2PIp23d/V3t22ZCWjPNVtqat+
ImpnzX6J4U49adzunTLo4N2bFVDlFBrtMlNVE2ck6+ye6M2DvnVk1Id81MWy/tqd
QTi3V8rQVfHQurpkDdt082FNnsTOh8H+CsfaG7I9rA5xaphix8nky/Hr/exkX/5l
LypOFzwRq8c8Z8xnpbKYWNUleNpPvYBLOgcBRoPAdr2QCHCJIodVaPWTZmqai2CV
6Oja+i2ndr1ytgq6is9gXKVqSDl9axHauoFdX/c9j/ol8A5cv/smqVhajHcGx9yl
yT9fwyk3Vf1uGLUvfzK/JVp4V6Vo93QlfleIvLU2HtsoKKZ1WGxSVs2NUtqWLmgM
SYXJRChgrnpO2Eu7qibhB7ZPa4bebj5H1TNx9axmXgiz0tGmh2iSkEvZEr+Tc84a
OA4QTk0jXn18KRxktWgp2LyM/y/b0szCeYsuP26dr3/ppSgOxLrHAW6s1EEZMret
0AWlgVw9lDrc+jexWdkRjVemAmvzeMnMLDDZMQeYj/C8I1L9ps/u3Bexb8YrLKCv
WtDLgf1kRW+8oV6wE7mDzlwIlLGWqac2psEXRzHTQxBA4NKQDKid+lQu5LN8YHw/
mBfLsucrzmamRkT4U1y5wSL16nR8NCN9YCsIRdnwB9mm/cNZiiqDtXm9H69Nga1P
kcMDPqR768LonBNOVo0POx6fwdtXMNIR3JdzvX2erLJ9VscfVtv9IjcW4Lua7Vvq
1EWKKQvg1w58cqNR1VrJfRmt0gzhVRwpozCtk6Gjv3M0iDY0USyMMg0jqXyBExUe
FobvWFw+rs0lOUIXT3SXOTY45I3sdnUKMnKCc9bEjkfB+T3Zorp2Ptlb3TiA++xm
0cpKZZlhCk+vP4CB2BvdX61ND4VKvIRLnpzgJCg7Du8wbCDPvvKTWUXLa3mR/nP3
zJf4KVXOYYN7uYMQuSVz1GP/xVo/w/x2JWY7zeF71AX2uZUDtkAoNAqCTW/UU10J
Z0CjcNsuuAMOjW/00nCECCrQxIllqT4WLbMKU4hpve4aCjG+5jaBT9eyeqAY04oU
bNqVK/tJuLPsdVozjUjpx+yEBgcLKyaoWPGUsLcRcl/dGHDfjES+HRPMThbnDvcV
/sEDydhbTrvxjQ9NIswn6trijJSsKcw0TmDCNTJ9fLYyeLbCH2PJRDCnkkVa0KV6
1eroRkckuqzT7BnSYZIdUHuePts5BYmKMWIW2RWaOHH16P8YQqRBAwkxqkUxg/bK
+OYVSEeCCuCCzTEVKWJ5hjHxsCj01Ivtbzr4b32M8SL6K/l/32QqDZokLkjZ1kvo
quvbeZzI861nE+W+xUlGTjEDkb9jUbCMUZz/jis3XUDDmZQRXAS7dOljYuLKRoLD
i8nkX0wlbspULvEEknbjYldpQdOzXa3QuapxeidY6C5VjiBkVEQuluTgayGyqPBK
CXXAbBoZ+uyL3tyOhiZ2AZt8thsjaQO4aGXV53EMaNZFwnSuHJGxwQwcPB3dWGjf
Ate2MzkLnXnCFnvIIt81yletk6gGgiWd7EDMLqZnzF8kpBbQ/+KtFjYXSKkWBm12
PlYwWFSCUhYLzHfnyQSgJyzeBhgKJiy9GF17dqMlmyRovR4dx/WvdqyNcQpzB417
jLK59883aB+qrl3zM2Ti1UF3Yrfzu+ZXvYEOm6MsQviEs6cc2PoOb4FjOD5P839B
6ca+6rXVyAHPdJUf9octWoedNeXueCQFns2DLoMq8F02UUCmo8JcE1sfjBiAANXM
kQwbbince11n7vKT6B4oh6ROblFBPwhXqaJpljty2jscVshYUSWT1Vx6FGQXAyNN
5AAejmJt772Gk0cJxMbR6Gg6PrHkaGiC1sHn7EcIW8EVPT+c/3MJgIT6SDXet7Vq
cuxzq5+szUwgvUEC4FKAhCBdbNXdXZaGudlRbNkWL0xh5vcwUYzgHvVjIbmGLuS2
9CabrXJLLJXTyJOrGnSj592VS5zJ/bGgEaEGHzHb4Tj/09GBJbeMhkEOm/5gsm8U
CPMNzJkmzK/KJqPdwGMxauPrGZCeseZ8d/Uz2rGCPlYkye4m5pRmBpbS3c1tHh7K
MEggcMdBSJN36M9xv0fc58nI3z5k4XKkFx62vvmpYneK8v09x4UWBXRInlaVa5M8
cs5ZOUy3+zh2ICN72GXA3yVwaANy//odamzGm4UYvOVzTl1arOwE8L7OF19CL7qR
pOJuYJuVMBsDzfpVQvmiOtML6YVMuXR0DIsbmE1lrEgLIuvzUGM4TS2jcZ1KQfGS
m2I0PwDmjH2wAw9+C+H1j9P1vD5JH6jMVhNlrcpwABJt1f1yuSiOoQyeTdopkckg
aum46I3hHXFtPCqnB2nUekaYNXjSYa4b/rY1X5/bt+N5+ixGMJUQtox8v4wt4zD5
O06jVszWj4xLHbXRaX32udK02GewDX4jGUW4ZIOR6nXNr2kFifjBJgxn/hUCilQD
y30gtDiu0l8CuFT8b3oDILVPAAluV9Z1rLdulBkbqcS4Z5Enkt2Yh9577WI8fxcs
HuzHWr55wJ6N/G/loxRoOxB2wbGOcAibPkhWle0uCphSE0FvLU2v5YlxvK3+2Fry
pmfCAPSoDbDH2zIAkP7XW7zzW8uS0iwFHVpMSuXS+ked50FIfV3I+yuOT/ixU3zN
78YbbsZTNquJKeD60ZNlX34Qw5cnO3EzHP2ugjeDgmipsHPfVNIHNYDEyojFo5B6
/h0JxHRLRtmGLtGL6TpVPTpnXHBSCef5tTI4lTz0qPUYGxiBHC7Z1xuYEYHrS+un
MWdWw8iaDSYEkpU2h2xZ0hr76GI8HL4mUu9+Hg02OLJnmgNTGLXORv1YIGkiPfHF
Qpq4n9zXy6x2tu5rmvhF7QIdP/LawEcZbER1GCe71eeCJEzcb7j4nsQQ5yyRVsZk
HQwijc/OZ7NCdfSkFHXJdW5GBDjbkR2fZxURZsSWnFRFRC0dQKMSrWAgxQdvqKHC
5Nsor7WYqRcRdyO2zrV7zQvuMZvoUHoidUu2tNUop8IkZ3u6vfAv2fQ98jBHvHLX
TL9eoGikzM+oRjJ/X44TAnEtmdaoKrq3ZC6Rq8pA+Tx7F/M7ID+m2Mnx7C6jd6wx
PrZ5RwBjqn5+dkFRokc8JJVgCQ/mvrRRMXYC6fEnxEoeTklZlvOwNfTcTiN0fb/q
y1r/uVdogIL1mfJL3kFULlyPygU1CSMbp7JB+ixrtfvgSnOu+0LfNORiS+PZ/qDX
u5VEkK8RLoZTUVqxUS8fPN4dnv6+fKay+KxEHQ/RQLiTCU65JevYXJcfyALGv3ix
I7ahtXdqrEqhMsb7atap4sCiKPEDJtUQyQ/W57WKJxAP5bc6c1oWssm6L1QutsOH
m/Suu5wfZn/5jsMMWyiteWEPOfDjaee1nL/f9iXgjWAZ5IA0boZFgeCW0CQ84VR7
jr49lob27jTd1evcwm5Bv0Juw+NyRokrgeTMdIPV0IL3DmcTK4MLmbEG6gZGMYuh
OunNaB4QfgkRkA3i+X298Nlh9MkAQuj6AwL15VYnqYrV8xi97AYuvDwB6YiUc/8y
VUrWqTpnJSabE5LFTsLtg4ujCEIsUaAWhwFAcip/u61Fcb91EjN0WWH9oy9ztw0x
hKI9aHfSfsFgcK2TLYx28I7iVeMA7F7F1fO/KWBVhqiSTLTU9LVnqaqjPEtEFJin
hfqt879iRl7VpzBt7xsq0P3uWGL+NMWsGKXSSvAU2sEPT2sfYt5e+9u1cCTteZUE
sOV9jxpp+n0/nij8JrS9Hhx/CFP7N8Gjc6AndRd/kEEjM9sEQOcfALyA//YRuEmJ
g1Ia5KD5iahukYsN2pwxJC3ArZNL8tMJzXFe/c9hk6a5MitZDL3xpxvYmsmgB1bt
6YeAzIYpFXQPVDhS3VIDKKz3M2MQXFX7hH/0r0lU+G68zscZf2yiH7UmxzdXNITl
0rOzOBjd4nAJ7k6RyTW74TcRfv9Q9b+0M3HIQlI+glZPMyZQ+9npqdA4J96reICe
Ho8wdqpQTgDJFx9zoOoQuT5aF7Q+uqX/N/qIFLWF4V7jwk2BByOW94RFyeQEGJeo
PhVUG0hFh1YMJ74gQW/f9GlQGEtrcJ35rnC5ttIFq8lGJTW3UXjpfOJSn9VPL4rD
9e72orTGSPjgCNuybLIG08hLVYzfcqWwfpXg7gR11gD6itcUmXyq8TdVgtp5K2ZP
Jzw2jamdpPPIsJUDyMHcjayTWdU1KGmcn6qR+ecPrMns9P8DuPRiqi7YyW8Fw+R3
StpV56/X3fVaoTkQ/+9vPW/r+197FzyURbByYResY9iElWwtiTJhOVTulfBDL9hu
bzcqnnqDeSKrCEHXz0XjH9tI1tQaYX8+iIBECmwWgWJL9epK8dojE8l2UWEn7CP8
cwHJCpGnblqk+iMxSW0PkVj+KJgbNh6dHppoU2y05mfQuzxLjShEoZMijO4nU3T9
PZTXJPvAiW7iQwP4ZazRO+EUTYn+je0G0MeasgP6X3mcb/Rj8j/Y+iLYSdfqfNEp
UnFt0zfjy1basJM84NcJgtcN9YEOOsOvI3fVyvcz7emw7EpB0OpOvMzwMzxc4JuF
g8vFa0BN8FKYET9BnjhxJg6XndliZzMh1Qb91Hgq05TV9RLUciGmRBtZzaSO8mPn
c3j4iS78wwbckKAQmydLqKMvcsycoynFOdDxUMnawBm9z/l7jfZ5CSSo5wqeUEWm
TX4MdL+CJnkrPCUf3eo3YJvtC/auy+rfexcLe6XQ4ZteCMdGkJydvTrDe0Fi3/Hu
gVgUPzdzea2J+p7s2lxxhySXqOGb1AfZG3HDr8826YzN1uARwL95kcWhSbVUZx3O
pFJdyC9ilsd0NMAZwhfrq++Gwb8/O73d/vhuFZi3qVdWkwiX/wzN329yaXRTNe+N
2w8ygvh2Y1ivKrQcoFPaYcc6+uzu36ZPqzkBxuTMkLP3sXDRRQwc9Samyclsaxrm
BWKvf++OZnun7E90Vvod2155hx64UKLuujqG3zf4Gf96ysUh34rcAfotFpUDH3BP
2/MvS0YxX+ckbdIh2rIQhumE9LkXcTdCrBqCOPWfsDaZ6xiP+8tTDW8SozelKZOS
cYce3i1lOtS1ChwG0h56Hp8K/PrMq+1WtvsaHquYeYXUxdov6quMIorxHHrg6tYG
/kcOPcK7tjOnF3s0c9+IjTaLph6+ghFDn5BU50mBRgbg0kbMSk9txfg6pM89wb1v
yIGaL0sby2uJJ8WxzS5gPF2DM6U0dvFq8hlUmIws5QfY77Do5zohM0uQ3+s5vJ/2
MGgQTmGu4UMHJ1W+7i50h1jVwDYrEH8jGSncKkrQxJalJwejO4qpaA6y6sAX3hWB
i1Bw8ngwPwpf4cYB2KKKqabo2kYyr+iy+p3LFBDSq81Pg0u1v/r8/AsUj+ovHyjp
ALScZRosEdXpeqNPLhSMRQSVGVyiiQMxyE1T6gO5JXbfMGRg5DnfF0P4f4M6YM/8
hIVFD3IKJ+SMBBLvhQAFRbScZNfk29wDJa2C+/5kqos/x0O8HvynxqsugFD7UbP5
EGz6P4/287gXWxNYhQA93PwDwUNajAfdc0JMRJvhNTMvK+FGDqAORS9vUT/k/4iq
iFmaTHUorcXW7Pcfxy98z3nL9tP95XBmVmnNHzimJN8o5CoDnEJlNI84TiTTy3rL
HlFNzWBJdtK6r8fvkn4Mw4ffgBn696Rtt/ojJxXdhFwNnPuoLP1VVKrnuJv7TJwj
p/uNSc+ri6c2TGicGX5x2BBcFw4xc/vfmPs/Ssl1PU8TgVyuFdp2dFmOWPeMmS+c
AfrCiokbCYYITt9hMj88EA1ZM3Xw3hyPlSR9lP2lu4pZnlp1YlEn02zpOXi4y4ce
7DNqBFvQRXnE1exmkUAfAeuBVPtPUVx6lKcnnkxrW5nIFWs/9JtNuOQ8/rpB66Xe
UymI0wxDODQr1hGFW/4+ghVBEW+deHWQ2l98iyXRqXJO12kwFHrtal3lbrKqjBbZ
TaRQOj8rw7ls6dINWTgHQMHSOoUsq3SpNk99YNxibSnoEInaesGvRYnDLEmWZB1/
AR9CIfz3awvnTCrqh/oDd7VxyDRZkOzbv+ag4KVu3VTTSNby9bO1xHO3VsFwPQU2
PMqS4srO8Tp+//IcBtjQeNi5Qmx0ued8GvSolB7ql6rRYJijSmycWYeZBiRUA9k9
NJY+rAr9ltzq+nrOx3eYX8Imt6kwIRmZVEANwQlTd+2Abk6fWwTKLqbM1Jngz4dI
wRRUkvhcABEleRL6sfkezZYj3+WV5WrWcAXUqhK2J65Ul5+z11nTgK87HkESw08G
N3GfRtyDxs9LLEkS8VDB25lKUB+9fSlD8qg4ESpqanKgdsTElxVZAGEqoAnM6pcO
L+sDKF4jz9ibHe8eWSbfGHNFDP9vzpRDKqY9Y2/6j69lSnJpsgg4iXM/lgwAUvPD
InCUNLSoRserNesq+BpWro/RaFNrhjnaluxAUHHaIJTwwEUr/DiXKAYzRdB+ug5k
YYBmBmftHfE8rXAF4e66knL7QUJ7ifWtXD8ARXYIUjrTgAJ8eo/RmNHU6ZbqoekA
54f4oLYbF2bqGllaeLfzzViG/EJTVo4k51LdI36c8MPwA4wsdlgSTge2nNrqSk2O
USYSfeN3MuIa+hYqlvDVLMtjyvoopGSSaXzkNY4oBrwAhQio/BEfXQHPPVHNC4YM
BV575RTDUxa+bQLmW4jhFcDb5WACFLz8/sBprccA1pTYvO0hqc68pIJKdx1Z591Q
AeDgPKvKp+dT6PQZWs5Pec6PaYUzG3vC3jiMKC5zVkihivqwQX6/UyuorbeGfQ/z
rGGAU7TMB6MBZ8TJf+3ig+WXPdW62CQMW+gkd5j8VC270lBk5ayPdb2Ik8bvS33g
O7cyvY3YjtAvGqnllZj2H8FwuXCx2yE9kbUlNe3z/L39VurglU+49M+Dv8wzqz0i
yL0UJ4k8mPTHj5+DcpOheribOlnP8I46ghIWEmYp++a+ZA/GO8opDmJahD9qOH7K
haJhhGjcLz8vdp7BkIoSLdzG0fsYk+tdrs8pv2Dzdn+uGPHN0t96i7/b0QDT9fuX
OelMuGbAFTHbx/uCj6/HkJ4sK+usIcCOjwt8mhzy2jEBU+8e35+1lrt7/bZBcZU5
2+WiAaSNvcKWihvYlrCTJ9fz5xNa1gDrsl14kBdbnMcug7S74PozZY7Oaf4DcfH5
d5rTJoN1vR2hOABpKbN0UeBe/zZGdDVITVXxsNyajxtjT4/a6/ZeQcbjQAPbyIBA
22eOZRH2G92iwDMgF4g2heAEmGq6qnHFsBhR6/KQ6ICBD5WWMLyz4n71nDxMmFDw
5IfwyCmWq87PpWT/VHYTuR1xdA7jf0cvgRZalKF2sp64TihxIpHnDwjojmIxS9r7
/iwBsioG/ZP2fViJP2IRSze0oct4Ui0SvBq4oSYcowV36qG7x4+OrS10tkGyN8T/
xGbtAZLQaLXgEsp6m/itXwFMOhzqLFWJ4bx7RVgjzz4zJQdVNyctht0b4/rL+o49
FzwtHHN60VsQ/IDg6jgsm4WxoFkwYhMIHPrjQft1W/E2EBkojr4FWVREcIRYJpto
x9e0+lrpxxnZWzuRCBlxmH7Ij8obo0FAKtfA0ktaZcGXDCVo8pq/a5AwHh23hq5b
D3CB/nGG7AeIZFb9iNcxbAaSbkrOBVvRF1Ikp1QGlYPgDBbsbhpmE6RojL9++Zim
Kef8b3N6In4OcpJ7Qghk1jDtSrnPldJYWBoQzqpY99ssNmAIrgQpahYVUSDqT0pp
0PBY13H2FBeV4vh/xBKF8WPkMvtITFgZ3jYCbOmQRNTfhLjAl6C4aazAsp/arkyo
DxQJo6FxvvcpewpmcqP8mHpZw3EhM5MDfAe9Av4WaDp+MGvJpM3d2B0Y02qN4Vsy
6hPwZFzItY/wQFxlj8x/qvRaIIUbsYT5iJn7AKNLjd3cBY70YZZOMZbUQJeG7au9
7wCMccJRcCYHYf1xQ5JUNX3XFL742lz/USKsBrQ8itv2ERzvvkVoKNZvYOfiSSmP
Nko65K4QaqOn+oZpbaWdfKsiE1IP8+KLc791tDvlNIPQ/tkeJhsbQy/Hexkez++E
//1djCiGUd/EkCi0OF7cKboZRgExwd/OLOUlS+njGp8Ur614flySo5KXojm/tHMb
V9WpKvVJV4GoCqcwnR64G6Pngd8ck8DcvHtagFO1ebj91gACTbJvoSFPGoHkvc6e
y8yQM6O2fOpP7QdEETgOWHUqxgUdKc5+2BX1FfyzaEFSv5Azqjxu2Ip9BVxytw+6
ysvvJzT26snLpUf71Hknz+v7GC1Z9dJ+PTCUlhPmK0KrX7OZoKqvdUf3kaNCyefi
/z2HJHKdsGmSVh20zJ+auPC+jXKzp8fL514nWcVI8bn/FI/5pMHw2rzVYNohRcwm
7zawSDTRLzEO2zENimHyzlrdWSkWf0f2lpDqq38GqLOPZ5zWo5UMuYe35UQAbkdG
gYvcHGnVhNpH0Pb8drkkIhoYpukZiwbtylW2fGcb+RKa0ao0dH+gyc+9m2i4gzGM
5zZtTEN3vnoFc+4s0MZI5LAfVGeKHhwSgqFbILMRSopKjPzb+GrGmMsk7VvCpxJo
VkS40No1nC16wIsoUAMCZQrJZtXA4sSjt9qJOHd1DlDXeFRVIOx2AoOsyb68kox0
0mgOONJDiGveb9PFGBbvK9yh+A25/rz7BJxtPtefNq1ZVZP2ABtTgj0uOoZTYKSk
Md4WASY3CptCvVyj1D7Qo+WUbaThPug4Z3VJk5H1wCJ1CVl3JovM+KSMSkDCCr4n
aM6fpMq9V95XtDokeeJGQDFhKiJJH14YLMOHbwVJ0ehr1gX+27iN36Dc1yi+/Pus
j+hQOgVwXYdLnBmr31mi3droRFPRnel3mNCq2+jsI9S2Oq7fJ0DIdWT4j/k/m4dh
o1/MuaYPndx2RoLAenyWlhtlWdJk6eE+ojXuHdxn5ZZo9+Z9/vNkMmSLPdA35fMR
5Z9rrwjuF1KyD5x0TffQAb3z1dj5UKvWzTwD1ocXuX/dw4ZXNx+4QcnovueZWrtg
ot5Zt5I9/oH+yVgzCkdcX/b2vzbtlDBAvqoR0nj7/3gIRfh/L61Lz4Q2AJV02Zl1
l3dAGaZujG24PFjp9b+z6ya9ha1Y5YU9CN4cJaJsvH7yOSMCoNugspTR2DbFwriN
3z8XE3oozKrPY+r92uBKJ8K/3J2WrSSP7RvMJoc6mg7fGIYyOTq33R9s/E9YsNT9
zseuMi6eKssLWdsDXDXMGYDAP/56hbZztEPqbWa8o6YqKmmYpVGjx+91eQkmb96l
/9/uNkoRizZ+f0YgYhr4HzC/J+wuuACGs53WciH0rP6OtOKreNqQ3y8K6efA5r9Z
NtGMgnt3eCo7W4/7XrnOXRyE0eNv8HFsmWnFv9UT/mhpTE8Pdt0IC0O/ABETHM1F
I+jcgSBgQGxQ3Qh+wyk6rlNgC6y08a0+N0yIdIMWFEaT7l1zfZWw7Mk4YSSxHYVY
WyqWy9PxYjfDymIAjHZm2RnATF8aH4k1NSUiimrEQAwoM53LCRHc9qnv2VzTQz6g
gEKNrbPbpBmBz6HIkQq3MnusHCPnbwqYwUfev0YTSZsBi5wfgt+z7/kOasXHAaRT
BYc7Zb5ErjwdzmQWaW8j15oPWI0te9qyhtD2plA2ICLPEjpwoC2t5oJmxA/2oNZD
1XNHvlfl4Q4f0X7uvxczTv2UhE4dgSV4duak1lRsqSoanjbOI2mFCF/ebjTRiBwC
LT9+czbIbkHYqfM90TvUhi5LIDKgRrkUjvUGrV81gPmCvZL+RQ8zYtXhIV3d13hS
6V6K6Sa0b16YAtluRP0tDPpb7OK0gsF7tYRZ4hjc9XfKwHHawHTsus6tN7vbVUEv
Wyj32Z1s8x1Bzb8DR5H4IKQ95TPONZY7wqO8hepEYr411mZXlEP1ubRNfcBmOl4W
oX1lzrMPCNji+pWz9XprIoSAY1SGXhMcudI4RYEsolizixS/4cpPU7MclB5KQcEl
cQp5LcwoUvY+YHbt/Xj8dGF3cgJ8JJQ1im9/I2lxinkcgMnoH6sDb4pbjbBg+xnG
J1t1awcoElFHnyCuV88/FPBmm1W4FnSfeI2fSDlN0XwfPuc3ruxCFAxplqr1wmJf
nMZy8QbbsOlExWpAOxeilf2fjV1Rioc02uHFersChqc4TpP1tUAqJVQ4Bt2+u5Nf
zk9Bg8GlYIqQBKl+d7n84iVhi7S3vl5JUgkYvrK5zpNV0dvrZPwpKBCJZsHM5Hmo
W1hWgHfPsHpszAzUoVCv8DrmLQ+Wcbqo14cgzMaJyesMBIETG2CrQD5cHZqm+Z1v
BFe6NRmAD96RBBhJIPpv9PvLhxfpd4vMBhEp9mE9ek7gyf4AQR4sk/PffXsxar1J
p1Wo24nW4yUwGhA+YfhGpNa+gEcB9y3M5R/wTwojBPulEaY9VVHg5yMoWN9gG8d+
IQis0d97virqAUf9HsMctUiBsJ7rjWwRx/dKQPf93sSUIWFkarNyJM4zZiZiRr6M
7bC0uGyIKgptyiZTUcqaH1UVqG/bboowT2ZbYEM11TNy6LLTH9nTtaXovBV6XgWs
5GlwruubNYiAbMebFz6Z/19wkYdRPY9C448+xM2NvvFaA5qXRa3uvweg7PsfzPLf
PoEngWXNbBgTK6yPsifippVDxtjO3TMWaVZnRpUx72T7v+tsX9E/F5u00+tE/t17
0taLcaeT60Xhi5J9JBnL1s15g6CN5mXgSwIHd8gw6IJju0IXXRzNrI1T5SEoPqFC
/Ny1u89MOhbbv7ZJu8myyVoc6wu2NT6KxDw3OPrpZ3hGYK1D9Kk/k124Oz14mtFp
CtvyNEKeAqLuesKOUDNyHwmdOlUgEH0DGOtCHCoIewyKWbmHgEIknl+kT/OTa4cn
HE4tl8ZHrSGl8PvYiJg1Wc0+B4xv4pD+Cq4cb8F2Hrj8Bn24IfWuKoL15BbX8Em0
S/9f1YXItB2xeHoFkn+m7QLMy+VQCan5HJMbnWhxeH9lMoj30kwNyurBC791eF87
ixC8+s1RVlnf0GlkqsBisRRKjAZggZyb4nzfE+QlKGMOcfYqj6Q/y/hoBdgcTXMM
ich+3e1Lq+TfXuuFLBCIgfQHdn1n2apg9o2Zj/yX9D/V+dJKYPU7QUQQ4eekmGtK
MUN63Y8aR8VyJGzPsp2OaRKLb7o/ToH5dsw6WQVAW84IXugsI20Ysg3JtQKFqtE/
c5f/StwR5GbNcLg7iWXMUrNQ8RbQigDg3RPJ7Jy1UNzio+7HHSGCzZ4lRlpUggSb
eQkYiJ/Tb9WGzLiHNQkXVHrfqAjWy5asqUdQIE1Ggbm1YwQy0hWu32C+Ab5K4UnV
iKEudYcM8vqs8zRQWcm99KzRJ7IAhVZHDxhHjvWSsGZq3feYslOWXnkTcuztMRuu
0Lw9Rn9QXuOdCHVRgL9f/JlIAQBBEru5REmtDHcnqOTJfM9sVCqKOpHjSI3flgWk
VhWj26TsfFC28I6R2xiUONJNwj2Ya+Lhcv2TM0Wgu72voMDnlomGpBeeaCRFWDtT
p/g08xPSHwKM+AwL9p/y9RqB1e2DE9CK0Q2MF17ljYocYCGq4pZAoJLJR7FylACY
DG4kr5KAxc9T78JD5YPU1o6YSxEj79FgjOX78KKP7keCAnWMyaKCbymmJ3zZzCMl
jw2bi4944sFlHw/DwoBusXUYwPHIl4qhdBfBj7oLow3GeeRscpyVkQe0dpBAq/+P
Ap7AB/ogmJmLyBNr1hyjMH2jF8NB/j0Yha+iDnNhDGEzUojMb0/mHnFAFSBvfIZW
VhSA1O9v6fYQZmm4+MmTvy9/cUm6xa1bil1EgUyw3bseWv3XkVkga2PbiH0TAOIj
rLJarSIvMP5YQhhIexyLCZ013SrmGfBZIUy/OKeJa5dgrAr45WEWjSlL7zXe/D6K
dlJ5b4j+kv+s+Mo3NVNWrEJIznCywTGGlVpNyqHCmQsuHTnOUVYF43Ta/b50JMTB
R7iuaAe1/S1JKcI3FppQuUpxQYTdI074optsYqE4mT2gIT3CGMPfr4YE6T/4jvgf
jf308uJ2798HmonuCBl8QtlOJeDWPxRO5HcAmp3tT8uhO8AXXme0UWajjQa5cq7g
2Vjv0vKi+EbTFm4km/a10g19rv5yUDSOY5IOLEdDOYP/nDHX9dR2oXR0QQIxUT4V
BhLzBsPru51aG6oHqke4k32sdF/MuuUy8K32ogz7MdBl8MEoiM74ysc/p6I19Z/k
NmDfv7q1VKAtQSZGjA/2JgWaiymXxqvq8G7210N/VUqt9wzpAsK7UT9De1RzVlGU
j7tvck9MM4mz9/qHaPAGgA35QABnHzoS/zIk49zk0O6n1nQHjQ/AKPR7PhlgFLUU
zwQAhIVrYoTieWA1jMuWl+LflzTylFprPFflO+M3XZXX+dQUBTWkEkxPusaAETwn
XkBKXY746fLXB47vV+J/mRUYDFzXqmnwDfHpN/XDSRPQyMe31xekyvaDRjchr7hR
GU/HSa/2MkzNXcWKtKz3p+1EbpQ5th57G+GVLzV6q6o3jCm7HRrlEjSfvuMKgT16
drXuas37mr/UKLpkCLEiKmDO9D7zbBmYDs1eJVt1hsG2g3mzLZDTD471V2fawWRm
c7iBdUwe/9Bz3gtky5z1G6ceQIl72EYh2XvDn6Atb+cinNgNLPNh+VLD31Ccp8Ds
g0Lp70uDX08IGPvG1fdZe7i5w9l8dC426EVt7GygwsPE4NrhreQmn6DwBiVgNNTb
fugIsEdxuXtdBcyv8LDuVweKYpCdbpiKoVs9eGqNC9CLeA74w0AObo+3KVBrw4Ao
iydDF+9kP58fK4Gq9RWOsZuV03rHRYXzbCNaZtlx8pNJaY/pb8Ho5XKz9AW4lPi+
u9PwzazNBlj33xumtngPTRAO7FAz9ghgiKsUYsil4NP6gmyo7XOKWYObV/9s1VZE
zDJ8FwL9XhNQXgZUQ1jp7qGNG4ATxhaDugFHVH/Ai7RNyxYRnAckHJWnp4laRXZF
6ZthfU9WArwYu+gxLCIGWgapuWoPnUItsGoNPKgejkBlO1WDXG9uNCxIb7LHK+Zm
jRkloVENc3c4l8y+SU7MZqJCVZKoo0gLYcyd5Xur5dRubFJIqqoEYiYLevugmf9x
z8uXCTZJmZ6fzQwPk1HAY/C2q0RVRz1h3AW5RJM5XVQfP8Lbqfy1ftqZ+P+qLZYN
fKowfwsX84FvTthzukODGyD/vyJC8HtpuW6PEoufd76+QOqPKk2lMYAT6Mq9zYa4
FzkB/hBQg7Kj2CeMz+eX6AmpslDiOgo+/VANuiv19zvlZw8OKAubIeZeRfgEpd/E
VM6GKwlvHYbSrCy+O3gllr5KiC9cnS+yJxJtAICKM8FJ9VNQMuDFppbakisHa8VR
GafNxSjvJRtK3v6nzF8EA8OaINpZpD8be+0QFH6t2HO4iEiFjgDPYyo0TY08JIJR
gM1n8p/K8R3wFpgrA9RNDkCZMu3pD1acSv8TQPGkTv58fCgn/3Sxk+/O+vbKkbPN
7AAZGy+IohxD0ohIW3OnsExD1LBaFU2BzZmij8GUzD0XWTJANnzHTiT9fFR+y8tO
Fmpkd3qx404K5ef60NBr2yiAKC0DJy1VjcQg8/eCClKd5AJr3q3XZcwyOW5n5Uf6
AcUTxroNHYlAQ3KNhV7123Yq4HVEzHRhcjjQ0Z0Lyp2HoOffGkQfDiWHU9uIQZLT
hL5SyX6zWyoR9eN6WspK2QHysIcTG5Fe3V3/19sacvO7Jexhf15mz+hRLKgy/BaW
qEupGZ+hSl+1L9QXQYGMD813yAhtuUP+vOJGRdGvw6sAJdpS/1uGjKp6C+qHeyom
afwGVFTj3KWn/bh8NNvYPUURUwA9F0fusBe0S2Q7IYq4Pkg5vJc8GCR8BrN0YU95
XV+gMyo7G9EMpnzcPEs8IadNS63THtpyD9VxIG6E1Q1FbMCpLDgGT8Lgm/8x7DkV
0pQ9iErQ8tDBJCAWbINB2TQ4haHPeD4iyO+96C9IhGo3x40xBzlZBRYoD49tF4So
+ikEfcfDVCzyWnqEMM8gABWZldNR32xGtbnFCtxNN/anb4tqSSiUErB2BW1MT2pW
0b3SJUosVgQS+Krh2gPnnxWv6GU0pRXFecN9wOi1g4bgo6c93msloyfArtxfSBix
+5ZwjkJanNez3E5u4WT4joXPhb/gWQHI6QI4PVFZ5B8z0yjYgkJOrIgWhu4EnvFy
UAT6w4/IEGPg6dSryfyq222/1SGCI+2/9M9cVl1u0nJUtkSe35t+mGktAGi2qorr
G3Qcbel3eypLTOcXJAY/gbakG3B3URJT8a7mpVbRHiYR1/m1uAmlvIWxevnZguja
yo949JfsLUTD0megRvTsqJO7iAxGgcYubW//e+QCkURi04fGBml4KJOEaxTwy6JW
9LcSdITmq6O7N4i4ELe9uqBaF4qhM5Jmr/fVJjsjR/jSaVSwD4M9lQc9P/jS+v92
+FzxtKSfaT6AvmCJPJ3vPELx01wfUxxrfBMooRKkqB1y3O9EiowR1r5d3Mz1Jean
/SoYOcKrkh+1L20GZOrkwm+nhtKzeqlQKGyamsvuM6LFRsefwnlLXRLdVqrmCsar
5GjQlkwpzbiJ9iMt/q+voOxQO9KzISbNqnSwTNBHSSD7zmCEkzDVf5Go9QNnk1J7
31yxALsZ0kz4GpplZyLLc/ER4kBWzivddMYMmDD0jEVZIpF40O1WV68o97pZp5V0
dmKZMmCV9QaM8CZL8KNTJp8Mz8i+DF/M+Rjg81x7ZnTPguJb8bPHUNiBVLqnuNxX
hdRdEH7Mjh2AxLcmD6j4rQg4a+/MlIn9pRnxg1ERbnj4sZKUHBTETB0tenXAam6T
nDEoGpbhUBpm48fLkzp6dXTZvvAUPaR8hi7LNEtat/D8s1o+fylWJdmJe9Wil/g+
J3/Wemm2KE+mU9Gk5+ybNOoMPR8YvNhiKx1jPxbpUgobwO/KUC6iJaMIZGWZt6zB
cZ1zIWAT2P/fs0cntzRGpPfOFD1T/HncWkdvtKmx+MqyTaRjB4DrDj22p0dChPfU
FoOThpb4bZP5l3mEyuHAc1DOEerFbHbSvzLwwZYB4Xm21VSmLGFig80FI8Tw1ATM
iu+JwHZ4si94rvk/ItZjAmLPUtJPalN/jLaevF01+OsNLKbWA2N85Ej50A0dA8fJ
Xe7ySDgSeLILXu9imcNqeEga/2fToUgJcd0hPxV+W/nbwnAZyEhhwlFsrLDSmuC5
oY3HX7xAz45ZAhqJTsymNSRr1uavNFwvvvcNhgLab4+qDHDyyL4xpTe/EI2uqhIB
me9QBR8/OTD4/bTnM957mrh3pNRqkLsvGkqDv8FkLHn3d4BbUQDBOJ/gWuhGzrSK
v0Rh8b7UVsx8Kh1Td5IJD8SLVmGpEin8gnp/BnFVLwgQ7/698Qgba3qIE1SVLSyi
lK4zrgOcx9r/RbnT0B7LGHtLGfSvSm3ZIaoPuIUQsv3iljhEOaH4WpawOQn2tVWR
I4GOfNJfr4lwmNG/+MjLDkdoof6ZJE5FjhtChGnTzmXNOXAer2Rwxmw0h3AL9Vz6
vRXSD58fzUHc22CLkHq48K7ZI2SjueSKq9bmn17gTO/Rto09/QDmpYTcDe2dYlkR
7uXIBotlST/R7dJPRQlAzHYMQFfYNbt8ChEKQwTOOlwXzdBCACV66HCciovDEesD
q/ARhUWqEFO6WKvtuLV/6VCEvCtmyx3f8UQI45s79Qm2LbrnkzSIJuOddVSxEilo
KAaqMmPmPLn3Aez2DQq9CjwBgBcYot34D4tYnhAviHRcn7RpoXt5oGwRVXwGnw9h
i3r9S4ioNORBVbqReqeHB2sCrJItqsQzBwnW5I8U3Rfc3jwqcwjHkXt/H2VzLbH7
AV5Wd2w6xIbQDlfgB7P296eCptOk6JYyjVsp1MFNqHSojtSrfErhQBULZG8U/MSz
qBTu7sva5dRHLAboFV983L+FScoc84JhQkCqkc2aZJrSLT5AdzFmAoA90V2/YVPf
U3ai2ncVekg0PFtjs3H+CvEQAuzSCyZczeb5QQbCRzn3AE+31JnYpbzPBLjdjnMF
0gopwYICnLDPxBrpO97dNZdYJJXHbHase6bjq52L5Gkvf8c7akniQe2S6/Y4jN4Z
qFumP6MNy8SbppmDeISMwmFXMV+9eKIC72+GkBuOyOWQL2HbrejYXmRiD5sISJXC
uz8xJuGFeJOCfufO0yBT84wgD7IpLT38hzDlfqEehNwsLpwcpdc9w2iXaRL1/af3
ikuIzG07hJDh30/foVE8BcoMXcqNCBn1b+P732jNSMKV8TVJ1+McCoAMNKLvg5Qu
xdLcJNk3qnZQ+B9Eo2vr5GgAb1x7LfcZQplrlrvNHRO3FXbujBccQv+orlXJ0ct3
iy8wC1B2nkoZB0cAmLhynhlI7z5NAqaoaRoxwJ20Fkzic05uZHgEZ345SXd7ywa6
8X/TLTtbmB/gafjWTwmG2ENoaGq64t6ps4MtHlIH8cxhHiIlKPwhk1jpMfYyfO7C
ej8DWnDM0iYl2cDD/PtVXfnt2OXT0eBKA8b+r0heq1ozDEml7QH1JdpgHVSz0auk
8S1579fxTr6BcNtvkfQX9m+WErjvEOpfKuO1TR3C+4jjPs1l+tS5piJ86sEgiZDA
EhOAARADv3dXDpFGj0RyzRTL5gGJG/5lqcsMlJy7JGaN8AGRIXBWVFp6KzGglBFK
cbT2nZFpvmTwA1dR+BjcTL0grXvHZwqSOrUvw59OkAfbrI5JGuOLx8X21PnyQzhs
DohQIG1sAnVlZWAStaej8hL7FPwGtSkbk8YeGoOIHJ27bpdWHbkZcvHwvI79Nmjb
6TpHR6mO7trITJxS/JwjG+ETNAVso6XaLYdeUZ0eEJDTmG2FIIO+jnv0PpOuae0Q
l4xH2ZSQmhoTVGLtK5yx7Jt8sZDlY4gamh9OXhlwqmB74eGpPKxBnl5calxrJDqC
ANZHe4dePS98gr8A2QV3CdQ9VuhAfxYPm7VkhIg+uAop5MrCudkroqbSj8rf66kZ
2QlKlwhwRzgO8GoNC79qYLRP3EP0SwQjv7X6pU04SewwCDZesTNwIHFMc3zYBgz7
lMloIJx50sla9RLm0xhfUV4T9dajmySTqMEQ62KuCSy2pHIwS/9yeHzC4vW/8GNZ
OyG++N6BrgbMd/vxl8MLa4hITml9NnJoCVKRK9soCOlGTWHS9vciCAV732d9zxUB
UKstHFsyS0SxSKIynkvDx/hxh4EHI61db7bdmUMf9LtO8Pm+wI+NFM3cOvz8O5Y1
bYCqRzjkA0j99J24HGTa50lMoQrEqUtE9SV9xAYPDXlNtwiX8zSxNvsnSjr4d1wV
VEpkmUj3PWU67/5cOcH9ri/zkZruSlhWyQAT8jUG4F5usAEW1A7DVnhM1Ixyw72C
PhzUZcv0+IqyyWIPRmoo2gyBlRhZyrSW7yiXSeOE1gQvyOcGaaJ/gbRRr6NmpNRA
nAXtoi+l+BkWrXgaKUJ696k7gpFofzaURXuuVYV81Cg92u7Oct/pXn+tu57hdsUN
ic4m1orxJF5Pd7aLuauEfgIZaeZq6qHAoQkSRX7ux0L5dO6tXmAkpfLuOH45GABS
KOdcMjaCsCRXuogq+w8caEaKQnS0dzv9fSXiBCfEFtU4W6EXN8Ayk4PHNJFhrEyQ
WAtlraZrDghS0O1IAbXNEf9y3J/YiXWORL3hG1cl1cMXRWSUuULc2QaN/IlTgFCi
OVkr8KEFx6lpw5mmKDXOq2DM73iK5e+CFMVIsFSFVDuBS8/QRZhoOAspeOI567Q4
4RVbjRzQZCbT32t3m9TKngh6hrZ7BSiDVxCPLpEpIPx6UEDRcWxW+0+hQitLDiPn
+2yrldopfUL8Gx0iZ9a+a+gNDmH1qa3A6dxXhoM92C7nn0rsVtCbuIdDRYb/lj0z
S/GvuyZblWJnkcDVLurDLfYCWUAI5aEymAzRVAZbtEPISRRwRYZNo5WLBVgTFsfw
ImY/iE4iNMGNW572OcUEYlQMxOCQMsA5j1ToZGu8XEqg1DRoXBK8IpRm0Da4xaUj
Z1WyvdXYH8Xbv6ovmgvXGF6VEgMuklh9N0SCCd8/XntqWlTdW5F/V5oxLbqMSrjy
yVUxlV/1m0/hh7wWrXBTGIofFw3f+KJOyEjz4hHwEi/F+IVpW37+ZP9n/zfZVBIY
gMDlpWgbgRvT6RvqlLEBsZtjhidJg+msdxrQzZ3TsQ/f0OZSAgn4cTu6lwjqFJnI
O95/HwO/MxwGP+nLAdSlebMkUx0b3jpLCYasu/qLrOlKTCqYnHmQbRPdaj8oPOhZ
ul+vy2C22celX2PGCDpJoHchlvewoBci6vTBbaNBn6B1OrBVGP9pNJqUTCKGD+sc
lTB3QfUysfqU5mvvqiK1BFscHmDLetNdkE2DjYW2iouax0tTz3V+ecKTjylVavuZ
LLfPDpgag0H+1O6WbuG80wRrpPN+bQKIANClPI3sIf3hP415NVJiAhE/iT+xW7ZU
J/ckSJkFpfsp/baAPcFKOYQ7EbUb/JNmznQNbpt8JDKEBA7PvDNP/P4DNhkbOUBb
1y0IaGG5bIC/dTBe4+R3IGs4FYZtc+SfE1Zp4MjaAzycnov6gOldlzaWujUJkhji
eqd+rheZvhNshvYTUaXY4TmS/nyLlUXtml1MTVoffP++JrkgWON2nyiRPOjdrbu0
4QalsIupW+5aL3VU4go/FrZGU9v0SiY8MDPET2jxncN09ZvFcAKQKkuRRkw0o1Cq
lLtavEqUFsdAlGNKxihu7i7MsNAFQx6sH+JDSFNzsem6qUQA8uYApMQ4DR4hjv5n
Ap3HyjYynQXY06JezdxgoecrxaiiJfXdaFc9hYwIbTLKi9dGFeqIUwhSfDfNbEMR
huRSuS21Ffcyh5ZXO5XfJA6UapySGkIdHHOO+GnZdjHxk6CjHMGamtsGcZPfPDBE
XTG4MpZpELRWzwEAjNvHhHAdq+OJ6fSc60UR5Za8cQi0K53bNSbxB/OtKQ8foiUZ
sT64fvPIxE1rF+nSNg+ErB3kGHQFLNJ7RmYKFzLhsyuq9gMQktY1U7mC4eD0z0Br
CZuOARCj72bqJZd6gLKgeZPy/QUhXZ+lL6kncX0S14fLBjNX5c+lLRPCadBtClZI
ccks4D8eO8h/hq4M5oCLv14hoKFgMHry97qtHatVHyBsn6aF3r7+ZcY1jp6Ve7+G
pVxWs3DF0zEevdNwmLgHt8+G4MV2EUd/L53TinlbWjVL8mtH7qfAmvmygEmF/fSR
63FwE1Bw7p1m9KMwX+BWoCaThVg3hNQIp40DXZO1ISTh4W1h0Yq6lVEY85ALCPZv
ueUY5owDZkh2kJUTjnC5bILDex3pb2wp4oNjmM9vO1XoyOZ9PeqASV/1caSajF0C
SoKlbYNWRMPdQJp/sitkcVjZP+PyUuEzAYLxw5GFUoybMSPquZXlF8qR+GbA9ypp
oHjbccfARNExSDti86X9ACLMc2x6f3JtR/UIOMn5HwCwXyl7rQVUn8mfj3npjvpy
QxNjtUDqsExdBsnYJKZYSxUzZ//ASDaCxy8xDrK+2kdyCarHmUnaMO8c3IVdtmxR
XPFcwhikBtY7+SVwbWHiVm2XCMu14QzxRIEZaaHecBi6gO56qyHV/Ba7lFTm41jM
r86CK4m5EofCtHh5eX/Cm4dLORFaA/aGqZf84VN2FGBjivEPxIbMbqXUiCkV2LaM
aGl+KI9X4tK2TOHOlauFMMV97ECH2ncemTDiHpU4vhCJf2nfafGpjzhRRbP1LvZk
noEqbehsHeBDdOU3AIrOMgbWMK2MnoatnL2O7atAC2juS7/b0irJQmLJWnu4uIhY
4j4y09of7fOx9DfzGYDGUk1/TARrdk61bwWk0Rc1afJwd0RzuafOxE2odN3YkGOo
FlJimJwavAoPhTJxNnuBUC0mzQG3hHzE3RGH+ixIhQL5ECtVo0SPz4sa9b0aBI3t
6OkmbRkEjAnba0z6/9p46mrISZFwUCGCHkEXXQoFhyXhSc6SzYSNu1/Pog70OxMn
9+t8HU6MFb0vTHURxCKlDf/vNYNckrKoUzIc6YVHmFjNTEL95sTedqTkjiNtDhLR
xcRh3Cfz2wYEKn8hUZfgJph1Mk44bmfIiGFqbvsSgEHF7zNT6gASN1Y4S5Nj6FZJ
qgFG7FeyuKeIH33D+xHks0FxMGC5e+qQ/5jEaafjtaxNZi4PwCpSAlMvIqP0yWwE
ZdiZzQtxUHHwUBmnVY5tEOjvh2y+1dbeWnldT+epW8VEvX23Zqbx7GMWKH6kq2rZ
EfPfBgmoQ1xp58MR2co9J1aBZYzlohYHNyXxqKNxMCO6/xnolxiuQGdGAlv+TtnV
WROIO8048Yn/QCCWAtbMdaZH+gxyERY5lPXF8mCCdQhaxt4lwTRT0CZPLFjNn3T6
2ajAYL+Hm7KNQz4r5C6uMYRf/26+Df0qigGVx23zucXcH7+FFcIjOczRfK9iTexE
0QErbEecQionp48xMjsEKdBZPbKgBV0qa9Hbxd56B+1q99RyUMv8+paUYJzrL//v
VcpJgfGVd4LPoScRA4bSpnQULAAz+d8mJix0GSQL7r82vjE4rEdtDDLe5v9XsFSm
uqoXjn1I1dMk0K1sbyEwy/PcGmJcpbx6+pMw34tbl9Mej1aMUSN+iTmkHTyw0vkA
4UB39PLd92LrdEPEEacpRqSgF/7shhPGUilaefi/hKvmGl2oURweYsQ5Y8tq1Yom
1tNRyuFLr7Hfaa8a5TK1qX/1UDny8PrcPu2YNU4SYw2k9s4B6e1AkZ1LUpSAHOUY
AR/6FTcZ71Hssdmwh5yKHiLIaVV1qqquuHQcYROgCKIfa268NWGh4ERU/FAuzgLz
oAZqI8NHsZO7IqhTz5pj+kloVkL0hk3i/TT1f6eA6LxkbUk6CtQiHNooCuwV05GK
EpOvcRfWKouT1XZT9K4E6wqEsGDJipV6/3G2O3xnq6kINGdGjaCKkHz3sL2+8SPH
LW75Kae6LB14j9XnP9ZQvoUoG+NfH3KoePKA0MKnK3sHIgG2HCm16PhddvtVvhro
+nTiPIvqzF1E+tPRFW3GZJ/vKa9YXySEC8tBQa96TMTbZGD2PWbifCWrUZqHqZ9I
IrOC+70XnOR4cc08SYAMmps67ZOFfYcY8cXQY8kyLbSHHQh7R/mBt1boE4bc139I
59Y/2ynqwMfeNaya0pQB6bJFzdA/fdE8YMkAdUzii8mv5We1xJkkRwWsKokLYPpj
spayb0eYgB4LiXI5IRdbNhAuGMhX+/Ozmft46/DAUMGnVngy5g6S3XKRaKx1SpTq
AdVIzR6P8O6DYcnaQxVyKUD9y0Args1aBvaUx5Ow3XznsCIvztKh5ooWgVmb3bSR
TnowtnENDVCYnNwsO6QgpXSHlJMyuwFhjurU23GZJmi/NpTojoHT4gPn3PE08yzy
/xW//TKyEs2YlMqNvj3DTN5v9LuX1oR9btHPzY+hXb9pA8FUWpksvD9CPVCnbysH
cunKGZhQpOCoG42P4cspGTbb+eaXDwfFNkkUrIBp3te8FQ3yO/pyERwTjVxjiDko
oGWI3DgGAp33Nrx0NmU8/aOnn7XV/ncbHSUBON6r6CNDwG3SeG5tRvh92JbSalSg
ClEgsBHKvGoF77SypHQgNa+4VOMiW8/raUZ11ILnBjvi89Xs2iqVDA4M2IGlcdZC
WUE9zu/j5HXPa9XcP10CUdQ8V6+97oF9PoM2T90dy62CAgDZrbBmUDXW3scT1saI
CKtxXEoOSFpu/0FZPtmkOXsVrAI8FBu/kT2K+OiymTO5xeVtgbpKUYd3WHYrrU+i
CuPnnS7pyBrdnXNCFDBeqUXKPEK2ds3Sf+aril0L97LsJV8CIlog1CWdIZUvCjvs
RuNPVDJP3qRT9FQd9F0+I57992v3TefK5jDDLzmuXgWW8+E+4fckOvvjcLYFbMzd
W8GBjU1u7/aXHLJ6Uyew2ArL4fpmgEmI81szs4DzK1xX2k5zdlfAh4INyrU3tEI5
iPiX6JjcBsvL3QNRrYZTN5J6vmxsvhmwWkDHW9sOg66mj2EDrHMnm9Q2nVR2dwzJ
eKP5Lvd8NLlYgIT45t+d2Eq64J7C+cD5rvJWvX9eNBz/IC4Jb/eCB3v5s/PHmfSg
8ULu8D5VW73ugnnX6sUoalnidOm/5Vctl3zqehx/TBZ6kX8TH1I0PsT6lsUq2WvC
kUO4eJLMwPF4srAyr0sRPBQm9wtvHR12/CMueCMqMYX12EgWH4jdI20PrSMChhtu
BVDtYP+Q8Exj7DhUWYYbVI7fqFiryXoSk3puPTSdNTz1zda/Rxfd9IVHWzDmYVuk
ObiX9mA94BvcsHOXw4tj/F3WnfYdLC9U4RWdLx383EDSPfLGqIf5hbVs3riep0bL
PxfoLVi08coDhqXaLvqAimD9dofihXgNlfaxhOp+jcFU8XRlwtGOitgaS2Bv8O0y
JHHMQFPVhdIfTDahXevMnr1857YwYuCFu/Ga9hRkYFAnhE+B4W/6NXz1xnB16w1v
lOPxe1HsfCJ8m0mZLPQKOuWHzS5KKZ6D0uNCpIrUwWdkfhaQTtZCuWCthVD4lbNr
C2z9or2ACQnRq3WhtVHrfGVRnt0/yAZAGcYEaotODyZvrGRR1NWywrj52NEy2Gjm
m2TyoxmHkUCWInaZFQvFO77SdepP4nmceSb4AMITMBTIg5JHFItfUOMNJ1UbPW8W
OKF14z+2ApuNO1zQzLEun2p8SCPeT7ANnUfME/sEmyZQruGYDV2v4ESY2MIE/WNg
HmuHWs04NhMgdgbTGDCJK5mURSWhqQ6S7Cq1+c4mCHnB2k8nB3zrnscv069eMK/7
Ifpno69SLspLvHOiCGW+pxl7KA5b/0kHFWYX/jTc9HXZhMvwyAiTcFgfgn7rN9Op
0jH7TqClRhjqC52Du+VbujCwlBkOt72bDr+bEACpkLZIV3BvnamEHmOcC4MYbH0k
L5QaL0MArkh498fzdhN4aF3ApiZ4r+Sy9RQzqo+2dSESIuFuIVS/85Rv0YWpSo1M
zmZPBw9iyok/RDQmWgNQnfNX2MuzMzg/+H0OFctceKXFoordWNqb2no7d2/XVTYU
wFEahI+P3CtbLsSFlNkR0kOcSXb1mmngf2mDzdZoqNpW3VCL9hHpccNPyrqs2YzH
inATJ6pZXT8URr7amNQJpArGe3igKrohnkXE/RXQm2vQ0mvlZOXxtZqlyfNMsdhs
SfH1X8nWmDbEmaYrv4bMCJso4DNdzLDYrR8EO5xXA+gSPYMEwsDbO0AJFyQRwTwj
mvgHS2AzI6ivwIkC/Gb5qdZcYEpKDzHL5pVlcscVG5Os+BMRKbnOXtvoyHhYfvsk
bKIm9ScvX1tNIiqmG1WCHQT4fzbfML90DvTHRDmtxOMyOZmg9Jyokdijdjov/yg+
zyVgIr7r1Zx3WaV1F1iHPaefCXx1Q9MnRJf3NLTx+egI5qTSIqK/ozIdRFd7Zaq3
+eD4RFcEUucIMu4ul4j7QBFXhiovPyi+k2gWPJBlvFdgni1JXept52x9PX5tgPCt
F6ctl1jE7nz8YZU+kqw7OA6lH1BWdSyMkVnCMD+0/7YLkN8403erkBk5z0sfOMLm
3ZItYH5o7zXPUGgoVCllSw6lRj04oUnZhrOHS8mWv53uRyKgBZwjFmXDvrvfY6b+
HO6VdVIEbGJnGi0nnQOVrP4d2FpIFvbr92BslCc0RC1niIenulNotPZ90Yq7S38c
3ZUH5W4lTMhc3baSS27dB9LkPfLPvmjjoZz+os7KbxbehhUitqSmppOOYpZp4HQl
VzhSojD+zd8RGEc7i3br843tzkUlWIg0D4RlsiBRsfgzKr6BUIn5LMYBQemdYT5L
Sa5yyzlv6N2l8XZvPiIHxEaZFmqVlV4x+OBjGBeBXhauWQQpWw+riOggESyHfsaJ
/+quNVzmvWry49iy0t7A3GinE83NrcWqTMTQ5nfdvCrQJhKpO1X5HLEDXZcxdzxU
glnTvRd8HXu5wJQSqLX5zQWXC1jdVexnz1KKQKUml+8H2bY4IYoLCwHadL4RgBo9
2L2WEhNy8SOcjzozqBQB3uOqWy2ch0+REqafHpEnOFHsRf8uBcUraCgMxhmF4I4J
TiFu88548QY7Nz1BkcLzmT7P6ISiHmdd4SnhvG5EX45WKv5Ryqev1S9Ktr/VfzDJ
++jrmYv2GlwrSGJ6ujH/Q3joiZBHG2/tX2VnYo9UjvOrF0eAVjfvQpLN/EcrJG2i
V2lwWshSBHtDPrbBB06e9EpiHcc1b1z7NDsYqLcpNYQQll3wUblfnQX0EA8GuxGJ
Fa9Hz75P8lAp6oDeGg68n5wV1CWnWHN2c0gwtrjoca3CEylvTZNXXthb0JO5aU+G
0tnc6fxVBnsEHHhxhnKq9SqNFnrJ94PqRB6XNdZJjuk56aSSTecfkPyfN7x4Lm04
vC5A//bM8pNNdi2jb7uF5L/5c4RoWQoBmjidKHdQnPJXldp+mr0N7l0kxKLtL2Lg
Eclr/OLWBrkrTkIRhcex+6DET5f4kXxg2xFCdGV7OpOcJt2+wd31a37uBvfirzXJ
hyK3OriMISAexMcn7xW4vXfYpxC0Ak2q2Znr7CAzUmDsTueD5i5gw+sipoxGjukM
+yLFgYI4Yf/zWap8tQUtkK2ZEyl47YM6ZeOZgwRmH6ylokem01Zur0DGMO+jASU7
2ksV/cOvoL2OJRcTbfRDWObpCIwtJcv0N9ZJtDvbkCEic9VWdp2wZ2vqSKjq1BbC
c5XwAyoutEyC9WaHC1NBNNzXONXP3Un0eMYsw+1lmjjGfBMC2Xy173nEbLjCydz1
gxNhcN3UAXol2ewGTZ3hw3yrzx7UZrvdRGVZ07NE661P+7r8pyeIYOt1vrIJ/ClR
6jPbVt8VVDLs9Nb7SVZzbdP+MieeClYVPcONHY8mFwqda2xqkJzfSzb4XQoJWATo
Qljf2HCDVJHJjqCHDwn1Tg2IkyEgZBX6wwxFLA6UVp8aMPfjhlc3vmfeby4H513A
hGVvQAim7H5Qks8wQNoBTYp/xhPcpttCy4FI4ZMu7OY03ERMLWmjYGNhswp1zcl5
QnX5VlM1iFflq844kjJN6viL4driVk3/15TqGNOSrk83yfNqBJ/b6U82quqspHTo
Kn76d4q0ktxc5mEz/qoZ0arG3rrJ+f4JWaJC44yx6zd+wiPTPfRZ9Ui+LCL5YeBx
7tt2DUHmCplBjJqTEY/Ci3ldzXSBb0HF88vk9ZQdxLpn29yNKffXDQDIJ/6JVFVN
GJbiTHOPK4MZSFqJpBy06358EMy7oUpVCsrFXPWTvC/UlV4t7J18RBtzS3yi2EUP
H6TPdfKzSgD8Twfz/iXS9eFgjBqiXlATHTf/bpA77gTCV0tU3azPTOJaQ7i3hMkT
kBGn0SsuXaxihJoxEbvqfbYOTUWrujorrTVAdbMnBQ2MRlYZh1BD2XcwuIVpqBhR
fYjCHBbeXLoHjuaidIpyDFBPC3ysghxzskMyDGViB2Ccg5S9O9YOdX+RWQufUHis
BD8jEDLNsCbPtKruVWySHyu5zhLUypzezDVj3aVQF+LSEB4UkLvI0rwSvGPGebvb
nPQxNWRXLXPFlOICcp0OIDW2aehi1cAzC91N3mkPbbWcYcyvlirbthJG2UBkygA2
aEf1WoyN/hzjdHBZ6ZHFYbCblAv2zX7lrO8Dm+8iyMAWLFzI3ISbd7/5hdxNDO+C
kaOT4JGjXUoyvUFxkxX6c5vUnemeJAAhsBjWgv0EwAloJkbChzuqWmELSPScraeR
hWMfQsgGxNLYfGJRCguk67Z6AJG1EBWWL4Wg6F3aR0IJE01IS+TcxmIPQYdwuKZf
9HHtLzjzvMENvw90PKa9A1d2UKIUrKmGh46kk/vbGMW3x0PRHWk/2b+f3NOPPd+M
FkM+ZwmqSo5FqMgC6xjoLQufStL0vDi+19ZgjPXUgIarQgOb8vc4W0syceStssXk
wzWzXZD+HFVXtvNIySw2HGwRd8hY4tVgjQ4mfBu6+gvOwngTWkOYgI3LbtoSxBdf
ukk1+2/fXDwvoKJ/d3eAj+eC5sI0DpSpIF4xLNtSK5Ni/S5QZAW8EkLfhv+3hM/u
6ec5oa7ry/26k978KLgaYV6ezNkkBba8U6a1OZ6Kb+6epGYUKkzm5Mkwc9vVLrEe
/5KgaPNxqlezfmt8DlNX6bRsDb1PnP3BQDev8dx3r69O9SX2YS6yzd0LB5XWxwIS
b3S6b6FxUynwEZB2fhQ3eZjailphLnQOwlhL9cPK09HssfOhrQkW6t01U+ei/day
mJmUVjJTpl54pzLddlXNe7u1iH7LNSoCuev8kHrImF5EgEFK35ChoGuGw9Jn52dz
V1uTVzkJG8iZyLyCrzwsHSrepQjARKcpWIvO2jCY8qo16PmKdUKRcrsE+uIIjAAt
kL2AcN2bbUaHfeA6CS2vCo75WDHr6aoSXl2ifqpcgi9EaYvqk4MNV8y6Kci0gakN
FHO0qlU/vbJZyke6NmaRZ7WUxpJmvVDv6Yruu1AsTibL5gqGF5g7B92UOmNNl7qe
QQ7ZXUszz8Zd0lM7OoQAATvGGqc4okzHk7Qrpgo5UnZA8F3ViFCOPNxKY6y8XHdo
tRCrs3LzObHHLzAIVD85ts4sd5kZn8Pan/mnf7dv27s0FWy0cDqt1KaYV6Or68nx
DI6NouvTT2Lv2Vlo0DFMWhiA6EXTJ5f5NZX+auBfi0rC/MBBgYbl+gs+9GX5ff7F
D06hqiagt/zGj7zUt2kBPovfRhW+haTfU5nse12V/bsPlZI9tLAWbO2KAB+fYcPu
rsPMgi7zC6oto4BFLliWEVvi3rb077pzWDAaWI6IKa8YuswdPGuXXT3IZ+psHHnP
vjpdOWTW5tYd3y/090WY1iercbAGXiLsgnqmauhSiKmg8RlHNpjNt1dLfQLwLJ+v
BkS3rRKYLTO8JQ8HMmK9sR4jTlAC9gac0XSV1RXwngLgcGbj7BCn0ufpIRmt5rMA
dsahZa7b0qy4GGTE+Jv59TljIWas6nmWgYuqWSiJZWx3Hg8w/rN8oTDp/b/W9tOl
a6XXJ7h5P4gaDwM0/FpU/npndhUXvAiCaKCv6gxPDckZxKLoTFOL14W7cIeffyOd
0csn52PDvE36eWclLnTwybexzGNuHPJniYU5d+071C4mKWzK4CsTDL59dacru+8c
vvXnDwHRKlxfwCOsbpwLsA3boYt7CuZTyWIvh439TpMCNAFgcvUGe6GotDDJ8PKk
A08SDiXbyuBOibE7D94dUOUUx8OuX/Y/LkYG7S7rhmooCEQe12LWkmwlrD5sXCaL
Sj1jGMdQOMAqqNryP86q+bGBVgEScbT9ZA1748iyGVkaA6TG8j2AhPjEhPCamb3M
2Rl8p68pkj9Z0c4y7s7UAi8J8RV5EFAz6lNDrhAk2nN1uGr09KK/UEhNQyqIsRE9
U0aaVFHtmAHWObFQNsb5B4bj+Njm8jeBHCmLiNC/TvcsSQIBMIkRv5n0uWkD4f0h
6qKRe8Oz4SLx8xeg2RMP0GjKN73VqwFWa+fxUTQGovtZbRzvUs1er6eSj/N74YUE
3Ml4gW12b1g2AHKK40xsMbIm29Auw1JpQvcd+E53OfYG0bM3+h0wgu+DJXqtzOI5
0AxvQ41fxcfmbB8f3HGUpFF5Pl1wb5RB6YUJGOwbnV0JkYrAY6Up551YT6zYlDPf
qjRl96iNlAXxXsYqk3U19Zcqk/9AdPuUdBOItAcXFVR8dlyQEMQ9lqIA1FqlmtWv
Pl0IvIy14H2zFNiw8/iV4twybwdu8rf3DI4Vt34Tjqm8aB63JL7MVlX3F+9pMLGn
L+9oz3CwFsI+tfU+jsdt7z9idtZ1twVkQa/2brIHEhXZweisPoVBCGwn6ygQ5qmm
UQd9ST4gFKxDOLR7sPOrEpm31LElzNMtNT0LlMQBFDDTTorjroNKIvRE/jGHoAOS
gLROv6aM2iuM/Dr2CvEeS/V5SehYCbwvdo9hWDJbMm5VPWMUcN2WmPYkXlCK5Bjo
x4ZbsB7433nDgr7XoGM6337CcGuf2xKOYWeXjWjv0kdm3UrTe9GtZuK1lHC9F9pp
3mOJZUCWQz/HkFpDkpAuCTV9xnCE9jafkjqrMrnv2OXbSSAjG6Nw9bEk9NnpZFBi
q1wSX5twVPvxqMyLyUCh2gZ2CjcCkbjH2MwTQOr+tBZPUrMUTdBZLPiXvVOKMs88
WRnf7z52jKf3wnYn5YkM5rP9amMgcDo1uxjELgMNXn9S7yBtpcOdnF5kPEToejj6
1R2KgqNOJ7wTKTtRghmv4CXC6vzPy51zYxh3EeZKFObKqpRIMQSM9olOg+974ZaF
iXm/8YWfeaedYLH7z1rqXtfJ4FMB6mHtQT2VHt0J8/VZWRv1552FQ0FqfsNlv6z+
veniuO4IpzOpi6zPqF6AZNgx7mtR8YHhgFNXrnB++161K/AmzSUPeyWTFKA+U13r
1UO/nGOLA4AR0ZuR5zL4uj26bM6LW164OMkIWqp5E5JZ0B1QN91aWB2tNM/bkRcp
LgTkmRhoTiGNHL3e8WKze8RBThssn4VHxZs+XnTJQoKEdwJl7bFoE8WCgJbs9JND
nOc+TFPeMgXyMGh5xPyZrkMYeHxsZxnpu9mc1ByLG75FzKHOfjRCrh6Oli+5MT8m
fcYHrUSuKm3JLqFmM+ULUrYQEzIiLJ+fxfijSsTru66TxxeOr99MaHk7dj+0ObaW
Vokt6yny/AASWfbUzFAAyqPHUyqb2czcPrWr4pIFsR0sEWRLQAQABE/yC6+DDPXv
FrijSAhGFrvB01ZrFmcHJtrxX2iE3xYWWBgJWdgbcBD/dfdkvnYrI+Zr4V86Xs9G
Uyp8b+8JxxmcaW2j0L04vY3tgBnKL9Rbd/Eb+/2KTdP9U0MchYd0bVXivO3CKqJU
YM0CWDitRN+Uc9It65QbnOquQ3+9cvgTumUFhNethOQE0J2dt+mQ5zYlG5lpK+na
dp89eE98UZKOpGjZ37Frh8dIjg9Wu3vNGth+uXxUygZCUpHFgc3TRn2kps168oIK
qp/Unkf+t4ytlyn/8OJ1ER0C2m5F5jhgy4fAKzjTY7dRDtTGVSDWZJpOdU8AGjjc
ZNPa6ML1NYYJT+tOKhHfqj7qzKxi9x3ZkdDGtUJ/28cyihPD2MznwfWFwQYBE+be
du5MLzvks/Hgp2+mJcgxNVANAz15lvIgd6R+EXyCIeeCYdX4mKw8C4KJReaDxpXk
SxToa0aZ65BXieodf6mFNUeEX3/5g32g/Wzpf0MijhUPSSJ725EtzcwnzYtG4xVS
aJH2P1dML6jHKxl3CBxsKWSznqw279+5OFDNbsuzcsni9eqUGmBFOrha/nLfESy0
spPR6ct98O6iM7/Z9VlPODioKyKRti0/JxdJyJFXIAwWRPeq0wIDc2iMZsBteDqq
LS+OTFh6plwQOiwugmTXB4wRCuaD5+f1O7SJmkp3CYz65/RtT4crYtoxpyhV/trN
Jfi8CP94eEbRepEks6u5h4igdDWmfYUUAj13CFf4tN2huXmITdL7ckIi+kxzcpgT
81c2Hpi43DmHprXYHCzrFKweTkeSCkMW2P77II9BLGGHRturHQgiWWVDWNHdZq+s
63c7HtvXYVF7sUYj9O5XqA428rcpSYFKocGh5BL4fTA0TZ5LT5Yw1gV1NEGF91z8
sBKIY/QJVuAgPN2Uefu97XQNPXTmtD0TAktMBA7vvZRvtGpJbS3oGQw6nub1mjbo
nqx8qPvrBx5Z3WKCtgrhD6PT2j/VrHb8fcXv7IFJyETQRWiifshjf1gVQBkl+JKp
sFVxsDIEqZPs3PrZ/2lexB9ePhAdV0WRK7NvHW089aA3fX8G81BUkAGRiAF+ax7F
3Lwv8GLkb7kb4FQW3qGD+F6hmfotDRYZ0xOl1AyLbmJCXxHkDU+HMiihwm2XK8B7
DPQ2b1mL9rZowjZvK9BSuTqWbvr7sVWFGgbcuhZaXiuHwwn1yOfcWChiwGUW2Rez
SrBQmdkrOiSaIn23w0cJT+TUQFxEIXvu1Ah2eXqaVODoiLo1r4p+4zT8f+XEyrcs
AIoCfK8LxJqwp2YZpgk/E3MoWJjhW78IwTd8kN4ZajZvNx0nS14NUrUv+zVEY0Oz
7AbKx3hhgIzH1/P4xrF3qRP9N6PiX7Z3kbnFX3pgEIcDt+xGEja/t7q8xvAgl7zF
9mLUi2Gayb6d/JFfS63Bth0xXxR8hCZHA/KB/LT3TvOW+5GH6t/+j64IsG6OsZ7P
mSW7nb44HvpWvzaGUAH99AvWGZEFLOTcXqYE4e0lYTVyWwZUXj9HuggGSyzQg0GA
YSaNZmfNQIBTGMD/3ICIyChzbOUoRy9X8KhLCg5Ml98RKZz9P2+1jnJ/EhzxSHUf
XUg7y7pILvn3a6kf7qPk9dqnq1ZllzPSyos1mY1XZxVPfimCPBPW8iNBZIGjS0VH
q31ql2PgcPPGAhzsl1EsT8QO7k+J7gLniD3AEcoGZSNHP1BX0ehkgbn8eRHNsImf
MfgkywXWB///bT6koElMCCXnO7w23xcFlsd2sLorJs7k4Kz0rQZCu3ymTR/SJs70
0uWZHm42fW49v5ccTHkYx+CwX7Vz0vPtynexyRf0o0yIRTsCpqlZfIdFtlGfv8Lt
TZKu04i5ylgAdxxxiShYpaoJ21CZEcMh8DTEbdLpB5opHXhaDjRbiewrg868iIF+
h9XNTuBZaiVmFIV6W3vwgm8Fi1esq0gN1dcU/g99Q8fIjHpNitp6kaEHiPeWpvQh
adbbLptJSEsS67dGURSOQQRuHShZwGO/Ht/aEzjJPJUqHMAHd1wfaDUfG5421Fsa
DJXfPd5/QQro228BBJE58t2HmVbz2OUOnRU9OGNTJ4hsCMBRk4ZWHxr1V0eaQlXa
3q6Jaxi4HlCdhdpiV7vCFmpBrVmWZcbWlmgVGjT/dkjfC+gMjtJxXV177qO/Q3MN
rRBXnygBlxmQ1SmLBJgLPAYnR/FMtCCuT23Ejkfo9XjzJA+BhqRgpogU0jnSwGgn
eIUtV0folIFtQmMaXhOwgpYwuB6NxgufGckjU03HWar5rZQ7/OWN023l6T2DNk3E
9KinxM/lZwiNUACxiPYiM1nZOadsgRNPLu3L0r+11HtmZiBbdsC33Nvc18gHtmGV
x74FoasBqpj11ynUYE2TFbeeL0oKhw0tENKN53kYgijTVWFVE1Yb11xXufSGyKgJ
9crc07LKx3cDe5XXnPw+b+jBg5lHqh1JmJUR9CxbIkJy8YCfxKCAiHnOxiL2jML5
sktQvRaRwHpugpSYgyizam7fbFEhvi0nO/CJ67rtZpu1zlk9zLbCDaYcOeWcocJO
8cAAOjoBT7kOwTyL22AyVFLK5m4w+qdfMzj6TM6sqpfPjxwsdcYs0mf05DlesCpD
GUIvZiL4zWhp/7GuedgOxdCaCqbf1Cddd+ClY8uwf9MZA4GwpY875V5TAWZt+4pF
for6Z82iqbaUJwkImWyxaRTk4WNCCVlnhcxgDrDSREopLGhnVRbP91s2NPDPFNC9
/KJopC+yehQEPbOs9bqquM8hVV5SyLWZ+oucS7WPOvIaaLEVQ53HOzCMUQ5ozfhR
icvtzece+pCiJaBcm9K2+eOZx9tfAeXm1NQ8dYNi9P6KHXI+77IxPVlTf7NhwqX1
IIYl1YuGrXcHW2udJ8q1xRhtgNu+ErXV468cBYxAS5CKAe6xMl/12p9JthH+8xWX
VUqAcpYM32lfRH7C9hU9VkNDVkGUqjXf4afqCccIkbpkvrBbt9UXldvv2HLvojSC
jw0Gz7mPmNZ61IfN+DxSSKhLp4krKyLq+VCXIc5YYZf8bgfdCOemIX41eeC/DNV1
Gi0Jo0uvxW3m5dL4BbQK5vQbBXMxvTznq24tNoSqzixQC4GDmebUhB81EqYtm7l8
n1gjoaXGDG0K0UhUtUnCcSZRD9vEnb+3aOU4RBVJzkQYPT7d9yphTPF3ky4VO+Cr
Kxrnlyvs+q09Pl6AygybUPACdvb7zAx9iErILlyP0i5ZCMGGZ+s8jjqlh2Kopp7j
B2uWs3FUGopQ2Lb4b02G4mLBqFobNNbebXWswKdBHsOzNjRd19UU9x+rNFPqrcqb
yT7QehhEfNV69XzV6OW7HkZg8diBrO/xk48cniX8YKWqmWx/juk4Mte2v0vMjliH
u2z+GSAmklepXlLS41tv4PtWhGRV5d7hJ8y5yyHjNCzcurjwRStD6a7Rkkh8ahNU
n9W+9qCM2qkVH3QLNOmoVedSaFKbN6l1LiKKw4MagBu391qi7mwBTinguOXblktJ
TjwhS7NWD36avXGqqtSk71qUBKsl+0LFuwdyMuTZmXdhjwKl65IAVNYGvDq/eZCY
WLG8f/pVBQSyxrYg8z6b3L3V1nLbKKBcQpX069n3xOTjIwPKebWZWpYrsD7R5mVZ
90C+av/rpNr7p9/IVaLXfZ6lsY0mP/m65eSD7ypQs218zC51LQhkUb7a7RtYbvu8
3IA/qFQc/bCCp/BXbTD7dJm+D2qyGini9alXekKu7PhRrk5eEXVCsL17PmZhb9tK
naZtMPY7Yp3PlHry3lOJKQcF8dEhcwr0x2F2CLwNOA5g5SPGEv8xKRXafbyblC5f
j1o3hghnu5MJRX6N2Q452X0WPe/k8kmDoLZvbXZNjcs70YrnjA3yaB+Htgr2CUSr
+MD6K7wtsoMMl7pgXWDpomamrf7tI6RjYReE8QATiPUSDoXHGK7v46OW/h3i6BIc
POzcUoFta4MfUm/mFfcMEKY0QSKMZDwQkrREwpZCpzlB6nqLkYXKKXm/4SVlwzpi
jiqYQLqed12CmR4qXdedbjdlg8MRCXDa8b22K9X7dMjHWmZPRviW40V4jZ5YpNj6
IXrI7H95A2vFzkCXZYQJ2EtEH6zag1x52LBx/cvF38LsiUAStxmYv7MOztmBcUnX
AuR1Nq3eC/7C/yopGM+0yUCQwAtBPCbgvuE6u+qOpm1IMy9hMYbxr0g3bYDyxSD7
ISCPmgVSulVyVF1AhpEuhNGH1jGv9jwRKz14wlIb5CwmugPn2kvp4r/bU70tbFPJ
hEIYuFSOyVmEFdsVl4qlMEssGCqGQK+5A8b8tHfa2cY5mbTKurEfE/iJDXS+ozqM
ZBHvmTahyUR6yUBLNpPWLwoCnRxDV87HP6BGoz+cbaqByzc44iCImMvFuQJXokYE
3Me4a1gPHR5/z6RjjbMcPoJYcinqtLR8RceuAyIXCa16ZwZVo6qlYQsDlQ4m1ec+
jhXIfc8uVr4uMTvmZzNiqwJjeBY0OPPFpqE4+/MHH7Qt/X6Sk7TPUQBdH3eaLczq
Qjyc3dvgGqx3Fq6598yrDTl0mog6HlHHGW/vU5uOWbTBge/Od77Nevl8BXkkg2aH
UgIHV8zOsfXXTx1GtxTco3hyU3PckznEzSn/ZmDiTdeB/OwNsV99N1aoiBs4cYrP
zweuo21rlOpumNTaN052UpG3bQMtnABGuTPEKpoNARpkOtXNg+xce8XOV31N/B3G
0shQwTWfshOzI8isGeUEDhFFj37RCzDspeJCz92eNQY5hQLm+Lp0Mq9qKe6YuEhi
UyTmSUjLKfoC5OdgK6AJkVHZk/4vxdyo25z3ZRwavuKxWMkYNrNf+XKsqJZmvyz2
pEyUK8KiaNJuF0TvVm9YPmXik32OcPiphS+SHz4yxkmq85n6QIbG2FVyrXdtpt1A
D5pMFdS4B4PzcUlbV7Z16fXb8hHvvIs6TrrnHB79eXAsDQv7kfFUIMT2jPA531kQ
2GcE6ApA0ZNDwARFcrOSIrNpbhni5KUAxCCFNTANGRG40h4FNZeKXLekyMbOIzB9
ZNz/bW9Wg0wH/aYTPvIfzd1e5x5tdM+Us8yMmzOo4NzH9RKcxyGwz1x0Dhoje4Gb
+bNNt4H2YEb/a8sZJt1jeXUV1AXK66qedMsrzc7xe2BmyE/5cIByZ2h/U95bkPeV
OazpKQDtg/laA8JjDjVRjo3g05gIkoUewRiQGj5XuNrVamkQTUr7zqMFMLKhaiAj
R5BaZYrwCTeTllRdXEqKFv0yrIXbnNexl/c5GyTQ4stZjNxQWs3vdlKSbC5uJ5Ir
hPr0Ya7N1VWEYQEk/VrIQk5ypEc0jfQXkL/86QDGS5oiePfzUeJMEm3J9fmmLcqw
YyRNhObo2wLTepEMelvXKM/sBhbqZIidEBhwj9MeydLW4K1pqJvJz3PR+51G/F3u
nrMszBJRRq4GBmp0E5eJYBADzTfsjty7QJavXawrw5/jEC1Nqs3Nbk7WrJXNICRu
7KJH7akiMtt8Z8SEooDoWcElMT5VhFI9YmMsGLeMMVFhlsTkhQE021sLz4zN1Ic1
SefwYIjDbmjtnysebi30EGAThF6cbCHa0py/sYU/4x4BpKp27ek6c07JKlm0aiFB
wDendNQgCfrll5+bnl22pM3SZgWU0MoECBU+CChcFC+G8fahzHPMynmCwjhp3PMT
9wVb+ImW2sQlpgNcA1Ph+Tgc3iO/lmJdwY+upLtGu7jKCGqjRGNOMKeV+P9rDEI3
DyK5fg9I9wP8UQtHR/CahhZk7B+owv9Qlsl2KjlVG6a67MRMmscZNEJWUFMZA/nH
VTRAHWPROqVAP67hvSFJvLWPKCDAD4ZhGkQhgJB8ETC2dqnLEFkWdOvxE70NNXrl
L62fQogZ2WGGCPyQ1cxHMSr5/jCdaHjCbOXHci2BSo08lG+gQ2LDKCDPwxixGAiD
36GgvGG7SraLtsvsYppopMRtbV4sbN2Zc2el1fwBqbrHuhSnJjZFCyyw/75gYPPe
8K67rXIHrcCnSbLnZ32Ihd5tX9G2Dlh9/otDF11C3w9SVGnSIqSeo8rkjGn01TCO
ia1oGCixCIqSvBS0c4Rhwa6O8pcnjmlY6G7RSHlnvEMhrkWVVDVGTGMODW12HtDO
ckC45Yb+jVxJC/MTWWvBkxfSMoOrWXi+6MJ0MzdVLSpYFrAXrJpa+SGqoBHJOoSK
DENlkazLxCNQKuIhq2glvMzwaPc3AD+7YncHK8i0SxvTKcH88i1kZI3PvaSFR9iI
bzxQ5dcPC3Ac+zqdM+P/rRE92T11XCQm2sD/SIGQWuleKdH7tooZitxsMBG5MlmO
YlM5EHZntpliYMilk3VZBC4Rf2ofJNPppnD76tcKwGxa2ZzQJjEDk46F1A3URWRR
njSLl8SNic9nW1h9XLEWwrzYbUMQmzk+RcPMEMHyDhf5RK35JQMDxqDxpr2Ib5sd
ubguFYIpJ8j6mxyNYXo2bF3OMwLand/ZQ25vvMQUPUuBW+aBLSrbD7GizZTQfsTu
AHS+zXv57Cr7FVzaJSHVDqRPLXW9ZxNAckVSJylwEeKxsy7jVqadF5v1xQs88LvA
GvyG6LvPcUCTPNKLq+NP2Bli3+zN+NxlyyFlELO1k60NnsM+490a/FD4ZPgzk2eu
DX7VAAQi5Sp0pZoVdl5RH7U6RMCxCuIJo66xMCkHFZ7FG+cllZriT+X54cxXIn1B
PJt9G0SC7B+zvXC2fhHXppfbMjdQsohVAkIxC/et4dSz9LkmJOYq/2aF+EawElIU
OYlM0F7gO8rBLkb+MpbSl45FXy0owCYFK3jlpo/SPLVisBeRDrH0Sxx5ByIoTOsn
HTd26JYf7eEcvqTaSrOsT8pTgbdxHBJ/5k4qRsas2NU1Zv4aThshJa8oTM0qw/5X
cqTW+E6g99lcK93s+d+1f/iwgRRdb6O+VortzyZdGQsC5w5eNgSmCWX0MetZJTsS
ymMfXBrTzhmP5AQ49hGMvYq9IiSHuT9i587FXcQqJaHQuxilb9yx5P4CHNj0m+pv
veh0rHG32fpCAXAdJKEUmdNJJeaCyJXYUFJXFHBDXZgaTCkpkx7fO77PDtDKNTgu
BcASl4lJkdj1Pz2eFJ+NyxWVUg6JcirqPhUBfs/ww8FQUbmdF0+1Ueb8h7xVGbMm
+kVaWynEcuPcxhF214gXuDzcNEiUZ3Nhm9oSUy3u61und1allaslX8gj2+xRhVpi
uoekF5vo+Mw4cAQaX/4s7B7ypuWvUKGJ4zvxXjA25araYsp/s4XDoFoUujFwPEjq
lFkHqz4O64UiUGwTJVF/DtsGXFt039nkO3RqPKR3A6DGjSx64O9DragIKay2zfp+
OMePVS70jwzUpqsBjErVY5jGOcLyP5UkNn7QYCfLXq+lRwAwyqXaIqNkeQzpqo81
tYMu837PN+fGsq2TIbeCa3eiLKnygkJZYVMUaM5Gc5lHowyMFMDOA20Pae3PLcRk
EMaQwz+Ebun95xg1Fr5oLRQTUGW37cuZv0LRJ5/o0A/r/Hk2uoAbUaDzfTarRovb
a4RxD5CoLnxbgDcHXg4watmRJ/0dpny/U+/FE5JWRRzeg8Iuh8l61D3ruEdMQUCA
mLr7JZ77Nf6msEI0UkqOmyqQUSzVQx3Gp5GjWo3oS0I8ZIE1gJizW0/Vz3BN1A+N
n6phsYGTIZcfoDWvAvO333O6DKRiXGEGnbZttwjNdvvw8cS85QV8bNzRobsPwAj4
7cD7Kkrjj4PhDDqokh4QW8N7KXxjm4uHxrIMJEzNTrOTrFXv4Hi/tEwU+usBz+Gl
6gWyVBxX5v8Tl/oKwgPBxsADetBy6c/UbSEVozQ68AJkaf6IwYmeB4VzY5rkPvpo
cbbLPlwG6+3eS6GdiVVjli2ngEWwNd2T0UD4Hjt5gij7Ssbjqz1/JBrRVmvHe77c
Tdid+HO4ALzCVgYwZUN2SFifXQT8Sv6PRyz64i5CFuljIWyjNlFwSEcOjbzddCrP
ycrDpxr6h79YEMqxeyosFOVFi4+TbULGi2M35+KhKSOkcPtFI7rGAz0nvuvL+hN7
HLy3P3v1NImMkIO8C8v/b0R5uZq+XgpLnbumdE8QnLbGdi9uQLIMpxUm26jZSyfa
wA6t38DspttLW+puJ7b+2JBSpl7eCXCNvhb9RU15wFiZpSe0e1wcr4YvM3u3eGSN
9ccEeTn2Ured3jruBn5oKS+MIW9E7VtEa/1uct+xxFGlzBjy3Do8HebE5iERFL/k
VjwjWA9VbgYoFY4PbUJtr2HCOkUsYW8Iipv0d1iM21aXsOHGaf8kaGPk4YS3F4t8
A8pni9K7RUYKc/d+9YS3ehnSljwjRkA9XjLE59IT15FzBYd9AClw9zFC7b2fMC0x
/k1jQZYaofGquFUR56tv7BcEkwdR+u0hz3XXAZx20ddwpEs6gBuO7mtFP362P8se
xiVCj3fYH66025hv2uCWdu2EOXtc+y271JFgYbNlApJJtD8aMPxBlpINdaySnepO
rumpwAB5dw2/WILI2Qd69s/mj1PkeX5s4hKGzIcoZjR10nLrCN5sKWO4KRGyT+Ti
20QLFP9NRkVWqTuqzDNKmWTQ0j7zDg/QUdqEjlUr5HsZudiNESu3BQR6U/WuX9Bc
6DMwY8y9PsR2ZuTNnLvY8zA2l7/CwFnrwqfX0cdv0LQLc4CJuSYFninUpDef94aK
QONFaa1yvPw5znBa1t9kFW82E5MOW40HIuV+ndwhltoTgwSb1jg2icUHZ//O0NUC
WIQ0NroBgsPWUNCuNvJluR0kdNbuEuXFNp/NggofaGXOVw/jbwEq4NZ0UCqwSiem
K4leXJ2KVFapUcz/3qlVOLDFT5ClRvhHvVAVeDercfhB69AMMrBB176vgNOempIu
RynmylcoA14y7BKMx/ObtlEGVEN7r+9PVP/NBY5ZiWF4G0XltVV0GO408PiqCdTM
sueCwLSzkYr9gnR+5UT1FlzBNxZN0yCAu+ZYD3870gsmSPqOuniRdKYOvxCAbneL
487ZH1nTDJ81P8RSVwpmKXWXCZuiQYE8lTxakVHS245EeOS/H40Q1u44WrbvdiIr
LXY4f45ePV3IFR5QWXqXbIrj5XzyAc0GHXMpDnsBxQCect152uz8GR+CCdHKIvBe
D19EynSNtEM6iQ4KFt8tTI/kI6vYlrDoEGEFtxy/a0JskYENHPtsG/ryXZFN53VK
+23T3H8qsUV5vPxbWuRKgIoudlMxW92/u4efN500sas/jKMjMUcrLpJmK4Q2dLeD
ToyLlliAD674HszlxbW79lAIqM81vpUXH1ok8yrdbz+spXVIy0tHjG7GQzV7vajz
uGQAmT0tL4BMfN9LSg66Ccs73bgcYAsq/A9ZrBZHln3DGFJv2YSdqSkvsMFchhAC
V9OmLqYx19jQstsz2srTzcCr4L1iNjq/qDBdNHzlcbshhzszMd+EK1+K2TWxsh/1
V0MgJui7AwvlfKCIY1IEWQFhYkP3vcPoAXEIZqzX3kgHhIZz7zxXWIqFbN+udnGe
BTS5Bvueo2gxbw8PIAFrGdUbfq0ioPph1le6U4IC4I1pNsskVl8RlPt6bEBup2Qz
F40HY6BYisltx0aaV02ABqKCZjuGFjh4MrSZinUzbIx/+fx4ucngN09DqCDeEHx4
AiCVGBj+4VUmHZ+0Ivly/NJh8uke62hSz1tQqR9CsjcWZ5KENSZajBvYRJrvAPVM
ba39e4qojKhwkPUeOOvogEqY+FRPHGua9M98SUgj0WdMyKNWznwBAx6HX/sV+6z1
SJ0ZruLit1gYNjHLbOQzwi7+1x7rIGIN42zg7E6AYLslegJ3APZPpNy3JEGR5bYv
xhs64DTWzrd/MUA7VkJuD2dtKfJIjK4GWalLKE8B2UXwjYPy2C7cPexnaOngk648
G0ceJSd4jS6wE/77vvLuniwlIiee/UJE/76omQ7VqQVm7RwwNaEmMNgfqKUVDpOn
s8BgwtNwbxIDabp+aIl+COx17OuIKkIE5Z8ht93g39M44igXHn1R53s556JrZBHC
pghaMnjQTWv6OSNMUBKi0P0UKKToVlDQ9ifJe1eTUYCNvRzwc68YVfBrIBhYNA39
L7auuKvT/+nrnc4pXBBIfquliRANenIQD3BbxkV4FBDXOYPh4CcDL++R4hrtb9iW
r6DK1ewKsY8OWon2W9saWhmNi5rxtkmL1bCJrT79kS6pQIrTwZf773A1W4JaqdVh
V4y0wq+GYsvqX9i4f9NVSPQWWOh1g12Gp+riaXeNG1JLEroiGWGvpHuduto5tUD8
HdnKY2I/2U2M5s9a1nTdeR4Tqmm9di/9jSQavZwWEeUbIwZP83Kg93duD03aQ5kh
1ACdzbEeun7tXg97KCEAzlrH1l6Iw/XpIf6tYkA2uuhVxusYuh+SIUw7ncAYdN/k
IasHZHDIxNOYogVZosEBRH+gvL9Ad28zMPHSPSIhqsBlFcih6ADwUS3lSoA2mwsA
czAFXuYX0jejfVSGUqab4yW2hCBPRhCY898BMjI/JOMPij7SlEcJ3TT3Jjp6k/og
yEk88mWjQCqrBjxBBfuJnNmor9RAXHq9y19wO0lyer1pDyKIdoLaY1fVoM6VNgUK
4oDlBIEVAlOEreZbDNMR/YfMoLFTkg9OZW1bGaNYpqKXi/OrBdgXVk5L/M+vdrZh
mb05MhCl8L/MMNRrNVXDPWS2mqUaPVOWSeYeqXgIFb+K18Rw3BOuliUqgch04hu+
1C9+cWTbK3jZwTkxbZ94SSF16qgFYrHOxWRMzVDkF0Q1LxR1argIGBlEfeRNRReI
9jYyaxNylpWR1jiMIqWOI7qZoyH+xmCcvpWrac0667oFZ5kbDsCLRwX34cAWIh5m
EJ7QU3zEP4FcJgX836UU6eERPVDQi4lE0E0JUKECQnk7hBgI8G3s5aw6+4QfWRCU
py8c4Xe0Aoi00PVM4vpB3ebgq2jy91T6QXKYigd4dHEoOOz9dY5wGs2KSSSsqImc
WjcUViOje8J3/DmQGGFxa6TqCymPIFTScMCzGZmjkuj85GSf00z7iGzxBCb7AbQD
YpgJnQS5Rb8E8heAid+qoNCJ4SAv7tbSkwmtYwzE1sIKWIOwVJNejnHGCPGyeHTL
ed1/Tfe/vM6fBZR++E5FboUtvu10rPE1NI4x018wnF5dgVb2CcEj2Uvronjj9SX/
vL1PDlLjgIpJq5MJswRfGm8/BJaEMknDw8BFuiuOcLEwvIgC9RvG0hHwTJpt3rKn
EH1Uo4lG9zwZzfNVM8fi26111F4c55ErLBPFvq+vr1wKaqWP+abGTCYUuMx5jDwv
dfBTvVU93X2/5Yw/EjOCyIgXDM+tKKV6RJMYGSn2LaHpeEOLfRUXc4ySz1VkJK0c
J0v4D2rYiGujtRGbxm0oi8zQRH4wo07TV0D2lmuQz1ZN6YAOS5bkoqlC5MpBI+14
+8N2hYRTXKY/3gUPuHZzGfTIUEp+BU4rHaxTDjgOpNL6+/dCBs8o7pAJeMMYcsB0
glnTbYm/VVS/QQvbODVW5KdGkFpeno2uXTKc0EuJ7SK99idE9emuOisXjosKswEU
fdhCYWIhJzMSyCRKgV0JYke35U2fMqhjHOQjRagtvNbKVE5OMLru7b5Wq4EPznHf
IYkaEipY/v7Xd4gz56oL68iwq149znPJritceKHO5gNoCNg5UJi8ykyo5aG5dDv9
iclS11xsbb7qjdhpnUGt8ZyAtiZJhtagr/2V74gBE1eNKVi85smX0MJ7OIehgzyC
zTNO8CduPoIAWLihG2RitHCciCqkaYoBdjUOPrvaNNUAQadndrjq93YM1j/QzcvW
dNP0sg8xya8DDE527OqIz/vQmHr6DHjp07tVxHu1y90yCn9GpvGnaSxn0KIp2qBV
REEApRqoZt2mWDN2uEtFYHnjSW5h0saItfI4gqCBb5jyLxAlPD/+AHEvSp8IZoW8
2oETMgiPJe6xcZw9ZMOrIXdrul4LWcEZFwyh6ubZTJiJ99OM6nMPcUAOHLQIpDkM
QeH9z+KogV+enxu2RypwABAq14Re7HC2uCFkTUoAYSVOqhewWtax7jgZ6qw40sed
WEPMrbRIR34eGflcBcp2JUiJJKSedXsTPUFFcf8gKHgqQEiEY/75F+Irrn4bxDlB
768mwA1EC4YJ4NHIl3/VNYE92tpD8knuGvdrYM4Id9kf1ddLKd82WcqP+Lc5kZlA
halTXHkKY9lUZ697tPRUhZQLNyAO6mTImvgMQZyqtr2wq+znLbYCqDc8VtaRPWxF
Uxr4d2ARDpeF9gaOprO7XyfwEzRHKCeeFE9+gGlaBfED/BerRW/ZO8HQAr0VNd7E
8V74QkUeAHkV58vdYjodV2X1kigSeiEB35T9Ochr56VaRD41D6s4I3cG4DcHlqOW
SuhBX+7MfNxxQq3iHweHyI0ntuL7iYh8+0Mj3AttCvWspBB8BLhf3qRzThnvT9P6
BKUHdnjBuocTMJ1xCk3S1p/9FJXEbiIu6bSGeovgwuAP8k+wvsGH97qbs/VEbLbS
/4Ez4h8NrSAMyy2LUDz6nRT/1eu1sOIUgsrL6b2IE846fkmGW/7TpBI87KHz4TTY
h9DbFpzJtMk495XSvqaxV6+6x5/ocqkRByMix7V9c8Iew1+5wltMEsPW47wXdIWa
nZrJxGcWYhk/N+9Sbg9Ab/kM659yzCuBLaL69mUxrD680jJpomsrOOQmBsoiFkkM
iudwTnm0bQgskTt6X9LWo8JHuILAELajcjkg2HFPuvgww7J6srqrkjqRUNr2j3NL
l9gKjOJ8JPmNNyQwA8hIRz5TwhFq6AY8HiW2+VUhnK2klhkY3hxUU+BMMKOP1Dlk
abKuwJj96AndX3WDB4fhCpO1U/tpLqOTAi5+bKKp07j0Zo8YeSYSVvlx7LHRP5wt
zai65knKaGHnpH4MUiN0eZMmA6VHuNFAHFHQIxKKiPSWV02bmMuUqvLkpua7MjAK
x6zmuqpszdKKNdWhAY6mEoFdazyHFJjGxNO+rQyrPZviWFhvus9modDUJMNAa3C7
rmRtajE1tkrpiy4uCqoo2VgDV8HYUrkwaxohMUcm/uBx0Lud/5+bYU64/zi4sqK7
wM8NG5cH73Tdsd4Fi2HSuhMcC7L0kLmo+Kr2ohzafqhhwifxNVGoQZXWh7wsn4sw
Hs3HaYcaieRRuJvN0LowQYzCvg8xixUx8qAeovd42eYPN5qovqlhrpC6qkzTsrDn
n6Z9z/iEbeXyYwBHPlecHFXPVeq5ACF8CMB3nOxGbV2gdHla4l8bFOJK87VVcf4/
7TKH9MKSvAiso8K2Gftog5ycrMbm/wod4/hDgYtNgVXV0GGNHcWSgyNQQcHzrzkZ
W1P9SDK+Ph4n5JPoZpWVE3rWn12f3/uQJ4d/sZ8kymJHHJLH3nU+zxQwsueMAX4+
mgDbHRMZUEXcc/2vQXptRXGWAVt6lMLRZesBZRjZHmlkPs/MA1GIwyPQ8bxKncX3
BUFzqtynT6Agn3S8YagzAyC90m7OPI6FW2VX/68cguddtuMMjQ4JRxwN1iWQkAOH
e7RPn7WoW74acqhuYXtPiEJxWEU63YgRqH0ZE1QKASaDTV4P3R9560N2ZPM86rbD
GW2uunc0h+or6Kbhmzgwu4wiJCFrxb9pVy769xpsG93EQfxwqvhaW1IMpWclQdaS
xeCYC/7BzH0GTBiXdX1lRcV9mQxwvqHfu07B7G+Uzij9PFYJIUBfdNL9emMtKMJQ
/Hqawk/RJ85fW0C4cJmE7vRCakqCvs844AuigKuFgr+7Q23OSIjyWP4FXOtNzM+e
4Gb/MPyTHi+8gn18LkLECBiwv/7Cix2FGy66JOflO2u8NfoexnuxwpjEljmTYx6k
WUqtt7U9t9nR6Jq1NiAgA+uU1tRbpyVDbvwz9CGBeAW7gJ1n8XDGwEF8ET+S55zN
m0wxJ7xR96C3dS9RWHIHOihd5AvcC++bHwT+yHG+ZSMxrvKghTa3q+h29bEeSVGN
tM7R3C5RacSKam5MsVcdwcuR4lfa1wvHl+dVeu4ufGVYmpQa3mvgXzetZ4UcqNA5
diV1KAVLtMZRUR6nqWpQ1diHcdGyVlpk6La7afBTjxJixS/2FOLjXTUvvqbiYCgN
PmC7NYJlQeHqo90K3SateTgZP0lEUPQ7nMB8uEs3sXKBmBgrfZC9IAin2sTaTmNa
31rfhGtEW8ySnOHZgiins6xqVTi4EOuD3gOzixLGe8vAfN+YSZHd5VvISwajrmR2
8+SKy88c+xyOONMWM0VeM+LFIrt4ou1QRPvDz5uxknKBhnWTdJd5L89ZNH0S+0H8
OHwi5yh4p5tP47ep2Ebj2z/W/kpBWI92yGQ665RFQHBpDlasL7Goa3NgkkzgR4j7
9+msFD8uApeXb+CYfBbnmIINwTsJfyzVHGaQzrKkEVxS2txt9soFh+LYtHUCExE4
BBztHoo5TsOzVvKaIGphmFZMGvB+KHAK9dqbwklBHf5CRQIL8pHb3kQGUSg9KYcf
9Mtngx/iaRg9rShOvTDzFEKv6d1AiCfvRE2Ll0ftwVV6iCgOVMwBRO97J5gCoyuF
5ZT1YD7RQ0cHw2chk/wgGAeLz+u8XralFCDDw22BK0sd7LMkUvQkY7Hb9B3bTNMg
f44QYmI3tNEc0MkxrbF4lk5jbl2b3O8LZvItUeejmzN8ubCYY9m4tMzJcX88Rehz
t4BsYVYZzXzlOQ0aymdlZvRw/m2LdW3EISKjw5spabTZLBHw80lahnB7lEFhzDPp
yOkv39zFb8wkT3J6zMWIKqMGgZc24k64Gjhu+rKsdsDhaBlsiBf76Pxcgo4sV0hH
1pT8jpd8w8PsuwEvbhBw1hf7CSdhssncs0C5wyZ2nHnZ5/HV5fdNHAO7XoDYOhYm
UCe+Q6ZuezE1nfdvGVpqmNHre/Y6zGTfYuVo8NpovQNlRwWJ4sS49PLeenfBFXJP
6GUw5VQ7mQDKs9DlPDtaWdc73d+b4VJpPTjh2oTPYj3ADOU8QQyKMFNMwn0MpPVu
Lt0700BUzeQc5riJqezb5CtNdvgEyQXpDfFW3NQBvIJvFDkDRxKAmKJjp4GzVssU
3iE8T5vZHejj8Dot0oswREFlYW3YtI/6jWvbp/P5jd33FbYRDC8FPpGaex/I92q/
r/kTmY3ee+Dk3VORwSriaN4O12s8wIkpIGNusvTbNNJMyqHw9vhAqA6R7xlMwxyF
OfsqsZdEoIZ1XMeLNg5hNLnIzR/8ssm6BsoZMk0JR3hjVDdr0ZQOXYj/Aekixzf9
3RDCiiAyqSbfgF8uUVUxy61oSLR/Ou43Day/WL5S3YWnT88YMD5hRqgBZJsvj5TJ
uamKDcaRcjWqzu8eS2cLtWmpsb07rnBJPKR3GK4WNO6z4gK3UlMdPMLKwCm3Q993
NoBnvp8otWQjgdYrDYkoJunINjYU0DIumKM8O3WM4pJEjqc9pqwR8k46Qx5lCPUB
eDQfuj9DAl2DfUmvGw50CujJSYJaEZPfzSKlPtf+oDZk2otb2NQJ6Tdi5C9cAOJ2
ixeaw3L9ws1rbDTtV29hyVk7JDuC64edX5kaKu2nqpWfYMsr9WmPPb8dV+NnelR0
GuBWGEZAk+hOL9tyvqHYzaVFZC4reWa/wvCDMRrhjvQ3yMJfKzo+JL0Lq1NKwmL+
Tk6wdG8Iw831ENHZMKmr9aaGRrzcZKOCkO5PEuKcMXVfW2VlRwbjeJPV/65fpUpX
iPvU64Z5To/HcJCpwd+yn7PWehh+HiuQ3arx4F2GMJFPwZnRKDUjh9VHFeYokpsD
tmXOWOnFdODXSm6fCieXIOkk45IND/6uemBPbphDpR1xiLZyBujjq/jWc/mUH9Td
1FFgq161JpjwfhP+dy2LvmpH/Hz4pQL5zu0AXdVT6L5/pCRbU/DapUSP8LK/6mJG
1fa03s2xob3h4ArV8l/rGl0XiF9WVFcL3lJd0WmdpRHewI7MX0Q8ZFz6ugMstpZn
uPkzsCz+myvVz2p+j02m7k7GjTt7YqYMPUgVy05kEbIODp9vhRii+zUwGavCAMTr
IxWmhjnTVVx4vq+pn3R2WSXfp6WShXdRliqVt69PJl6ZN4cQMpQ0u4JWe2HbJGJD
xNCcAdxRyUpu/PqU+lNpc3NdRmHTdOb8UlMJWA+9Jv8fZpMHHn+tFz6Xt6pdNjBb
ykgLvyQaLK258nT/9lTPzKkv7PyAiiz3aNXqiBFO2RMx8S5gxI7fPSt6uJrvrp7m
fhkZnDk1w005UGg11PnqwtYO9QN0ImmkwZydPboSgSNWkN921ie2El7d2HIFC4IT
WPXuPhAWI854xn9ktwxYI1O74e3gSBSa6FpR4pGgI8AXCFR6G/whRBfqwUj9U2je
oEzAJcuctNYmkT0BUtET0rb1IKCfVrs2IGfhvWFecIXb67x/ch/oDyuUZIbSXzpD
RiGek4LJfjQqLyes3UOC33V0SawtbGRVgTdR4ED6rxPm+jD7gv5i5Gy50Be8zDwq
DjMYxzmxiGlqMnb5ciKCsHq+7+8XfrIzF1+RnVWI2f2abABmaHF3usb7EJYB2mOu
8ms1NaeAHKCy0OBWoM3MGBMIX1SjaR9uOprMqLt3FFNKQJkS+2ztM0RVfHK78YVq
ii7+Y/AyQGGt/j/UpWXsN6d8Flm0QgjvdbgbxayDQ/LTUUOv2ZidgvXAA4Mo5v2r
8xakMWxVuJLSE8ImBC3RWD8Ry3hUqTSm0kqPsqzDdtH2c88R9JgwltcUI4cO79j/
2wukYtaUQThs0NwTCVgD3teJ9cF9nWodcYHnhjW31VAKqjicL3JUc1qM8wTUKSkF
KuxqYVMlrMgLvJFGRpQ5POsJ15N7qYbqnxxd7UoruCpYYskwHs2dxQ5zvGBtFmrL
MKQHjRKS6U83potFL6wb5WW3hxs8cRKBAuNWxDQN83e/IV1SzxgE4bwmGKQTb80T
nuwjnguiZ6zQbj927U61yKggeE62fBSFFQlXSOvpgC7aSKFTOtlOnEoc8VXXgcMv
hfcwupMWmU/euemGPE7kHYhaCuSVm5wfBOxzv0AQTjA7zNgBdH+qurjC1TuCiFPo
RgzHJHeKfjSE8ivakRZTpiLpCfNHMujrEaOrPvNUqcchLPHEWp2KKFCl2dpJzk+Q
cNOoeEfvk0s7LQmeHtMQ2TcYJnrIvBukXyCJ7j+ZVQ11+Y319fZMBRNjViYjzUzU
Lgj+RVEghZZMaSto1NmvJI0AciqAFD736XHNo8nHiCFoEJAvRxlLlMfNGS21HKiE
YIYSugWFbTmTk0BcaVN617GLgBlFZLtIyC40TubMvhYZUAi/A38aMDMFnm6m6D/k
4eMc9P7oeY9BDq4luuwD5oTxrRxSpj5hbkO0BLlhsq85svRd9xtHdm98xwERQ1CF
oXbcZCZimprlTsnibpXu0dcvV4JM+KhNrfnJ9k0PRujGG1c4b42cvBTtwp0Hl7jf
00ED6i8xrvJEJPpzVut11mTbWn36fyGCFd2wasdOEwQbxIt3YQwmR10Z9KQcdQGA
Q/k8Hss0uqR8mAyDad1yTW9wUAPwhapo1yuODxqaiQblrpbLVz+W4YmNcgtqMkkR
h7b0ky2gcTBffbFBF3EsCPQL+Z6vAtcSOtbKhElHdf2mnpf1Y9uMHcPCQBz7Cw+R
56s9kacDzV8TkIl/d8++9fLN5lpKiejKaRNCL1XoR3X5W+6Jtz1VHreIcXtJi+kZ
c8K1NRm2GK9tKuSapVnSHfFgvVFFYkTqcMQtsfl34KFu9x0hYcqeIyearWIrhjbC
05qyOvRxInN4JHo/X+n5fi9cfV61b9TNYPyF9nwARsNwHid6VJAQvvCUwU1B8ng5
Fb7xPswBduv0MXUL/ccsg6QL9emdZadPSA1RRxqSXQQltIYSyGTth13ktCuqDlfa
DMHpe/Inu8hLcf/fzuKbFwlw7Cy7/qJOuBGfDLTfKE5W+VNhrkjce7oPtF4Dipn1
NxnaV3oUtkE6VZYq8lm91RWxuc7arJfbpmLP9LShBhyUDgCvCUNRZckPJiMFj7XV
pRklJRF6LOYrnCdBG+/YAuJuzq8ODM2mxciRKyKX24qfFEFiWsnaxGTm347ZPPsE
fojkVYDB+Zr9xLqMRVsoNbJO2OJSaIRvYQerbyA0rgV1r4ZRLzN72WhengnQmPiT
r7bo93zp/QNOTH1CTk5N+SluTbAx/MbxhPpBcrM9qFd/pWrPu331noNN4pSaa2Rc
tXJ01c8gnBrP0FK0OK0ugInSyyWo2R+Hdp+P6bzSIY0Onzw+gU7LaznyBg8TRK3/
/v9rqyo/6RB6H8LKqR/uUPpAnGoD5b9LyEMpfsW0b7iDz88rzqZiI/LghSU1F8q1
StksHS1UZ7cYFBwwMi4riCAXgaIWj1wgsdjpINP16zPNx4z6Po1N2OxLyYdpO7Tj
H0dXwAEpEVOpr9XFe4CuwCMAGIuKNWaDlKkb0/T/+RUr2dKluqG/OWXJjG8EAVAn
v6e9H4dgve0gpdzqI9y2sn7ZwQ5tYPj9yW9VmpU7KbziCkMa+6Y58ajk98w+sJyd
bjanrOxr+FjSsPIunyNJTAzlu7QO2BPG60kMZXBrOJXRys6GxTwsossN/bFfGmEw
+41zuYV42UspJjgeEewCLzLOGuZHBcR9P/mswVJLNROsKsLq3LY95nNXzmK9/0Gr
sjBzq0lazluDEwTaNmHH9lN+FNxQNJMOsedEx4I0Fi0DXNebGhjHX/jVs5CsYBVD
gtNLSFvRgx6uwb5cMaS1yDPSnxnBBy3mRHT93CIxROHw5QmxUjG8FbilDKBI01L4
2RDwwjwdK9jn1kVX1CoIvYrMgNxECJGWTKS8IhOTVy6nkRrK3p/kgT24pDms+yFJ
rBHYUvZK8w+myEVBHTE4UeSTlLX1Fyg76/lMY7O4QEzLc13UI5qdYgZKQr0LRqte
i4KGZ5A/gW701bNxHh2paZn6MLCCXknCdfNZ9GT/faV0e3WqK2g9xtvb5vP/HlJV
NHBzQvBCNCoBrZvPcSxYMqe2U+B0+VTCjV3cOCp34SsDbfpSdSfeh7Wzra2Ppx51
VkE6ujxZ0h1Wek8n/7tR10RzuzBzl7QBSue3YLQSRvYcTdgrMxGyMC9QhDnxlMpz
Ain35+H2ReA1UbQwxY7brKbY12ZOFaQ0xMP/WRXo1U82jcySY0qDoVCYMRf2NDkB
0rni9NlqVywmaIic64iPtAHOSIOztOaz59R++6WhuIdPtD3NDuHeKYU1QZfvFwbx
yW3Zar8+iCspBawPfFdkOhg6kduYetgj74LbWPqynnrBGYui7SZ/GsyfdcbLESuD
IwzSQhf4Bp+XdBkadzJAQUW9OuihSs5DdtnUz8xWO6yWtGdyyVeg6ErDRUmTMruO
Vaa4bsTgBWkuAzyVeKyIrJZ8Hal5tAfnjLmGWxpqx8mVGfYKaTyxEcoUcNFzEL24
owN2DB0f9A5SZ85bbpSUX5DTIk7cF86dMgomHrHe+lMIhX8WzrvoQ+x8JSrNbzgf
8ieurjB9nY/m3cQdQCFfX7ZsjyBkdGA/g2aw5Xas+dUKbjTovGWjlI+q7/hBYGxW
izyCG40e84iImvKBVCQJ/tFHNcppNnxu/Igf2V+YX1cYZ62Voqjx33SGy033n6pL
7D8qwX0Dg/+1ctISIWshVDGzCYNV7bIj7WPgbq4v6fGgbCy49PQYK2R04E6lBc4N
+gOordXKvEFb/pBVM+o10RkcqJFzZPz593fMg9fkUE1LIoikzS6kEk23hk2rfiNP
5Mv4Wc5M7umiZF0vC3yj+u4cClQ0Y3xp8PuBJyGXq0ZFpvn5gWcg4kkNnvB43cVW
hfw+Sj/98XsKkE6RV/rFvI3dUytbHQbMiptVSzgs6K6Sgax4XrtQ65OvkDOllKvY
AnqiKOOpHzFlKAzBI5DSMtpgckqp7sgqxd+Tyy0EwbvZwnBTSFy4CkqXujy2rtmC
/BcTk/678fzNSU5uvuh1bpj8+xVffoxxBt5o6B1v+u0GXnUeoJuqC6DyvWlPLtmw
8P/aLIUCGn9p6mrmyooHklC1AotSMnLDJ7xNBPnqRNTPLuBuy2UZKdwN7Cm90hF/
cDDikI/54+vshvT9fFcVn3Pn1K2BQbXjmazCzddYs2WBKyv5MIj7bokV/e37a9yn
860W/DavPta/YZRgwPoQ+XjwXGwuTROHJYOOeshos6LgyzxjaMH/hudGpG1HOEB2
9j2ohBwqJwb91XIxgALZhLMXp6KGNw4XdPgNZY+lakDK7lk6eGf48Hj01jX7G9nl
TWS6amM2WI/SgaFmjZ0OJ/oovip9gl7DYgHBdxg86xIJpSa/MOV9vrSYZ7+yBbsc
WihhosKKqZRf0EcoqPtmEocTPYTonAaKvIGUYthlKfSboBJdg09YFrFhv7fv7Qw7
6NxEVBAbq1+GFf4UMROHscRze1tKn1MXG9R1kTL+DTvjpFFF7ifp+gCjzmytOSgY
KVx/1TATDz1Q7PL+lbrYkJfOO6VKewctS5fggJzDlfxP/CH8z1PuidFIlPMaKsaP
RMh0tMPFlanDfCslpx5KAnk7VA/TJS8UFkoOWLzS/L6GBtzu6ml6Nm6VeiDy97v8
y+PLxwXFFCVf9sB38/rmg23HpVYLB85gVLPw3FhzhNRy9V8YUQG60RrzoSlWS4Jm
dRErich94CQgdX/QJlKVzVmQKrTSaaU4MwybX4PveDG/4JRPyk0wQfr/5ZPoSBKr
THS2SJW2eEyXffcKmm0pZ7VestucrZKeatdigty6iSPaLuZ+boxjEc9YDZIXaQqn
zIVkrQpaBJvm4HJ74aWLjcc/Cezc86wSOnyGjNmqwWMSFdKb+WDjw4pmsFQJaLZC
tOQhbXjyfJkPnuURC6dcDdF8aqNmQGfwOE4FOabBQrmSdaBTKQcmyQei1lz6r9L2
jAHfxjGPp+V+hHQhHgAdA0dcb6pHsiqrkMm9mXRCCxHriz+BUaBMwhMf+0/Yl88q
/TB5Y8GEKC29SH+2DsudZHYPgs7vmecDEoO+BQymzPIQ5a1vCH+cDTHeTtE6yzK2
fQ2XO3N5BaRcSstTJconm7+7tR42QWQWU5ophG9Z/cdK7DoxZ9NPwkq10CGgAH0y
Xf2dgfqcIbxWNO2/lB7S8gia+vzDm3gSFQcT8715iHZBjZl+UFkhVDMg1hm7u7Jg
2fmqyRkCYtncvYOKhJv1saCeMNxIBVHNfhA/SYNaUJ+/GUmMWf8QetoZTunKLLXC
OS0+W+sKe051cpBub4m3UfGCjSRM5RPdt+nglvg5e/hxlfrHV8OdWZxU/FumhDPA
uHx9urY4ojPL+kWClC1jSGO3ynxbeZRF1Zp3m+8veXiStWm8Rw4Vy8jCFtPGP1Sl
J8/uJXn4rhBWTCGfWmwllXIIZETprMUcITt/kcF59FZZaFGpyJL9k6avDCI2oSGs
Lk/1BO/P36+xogFxby3/gB5CBP5WoWlZ+9E+hO/Zja2YdnAEjjGopA3rvExf8uvu
4+nL7JczoKLBzT++hogeBF7WaS6xXPAK65Z2xOfmnlap6FmQm5Y1wP9o7icR90dQ
y4MTSPsgX79XIZVA0aqJ7f9nvc/vGO6VNXtcBT+ENYJTqcnhILeQIC3yZavAd/uQ
NcR7DpwOtx/ew0TdC3c1ZjRYkH5LzkaqgERJAgM9/ebofgLzvk1YHJOyNdazQtEU
z/6fzGX3/FNfFiyxlbl851Dpnd+3Y+xzjzdMcqGhvyAiKhyxqFHPJht93NwNQ/+s
mEGf3bpNxDDWPIuKVuTq/Za9QPk/T66AWvQTWSrvZ7HgbfjtWjJjBgu8Rz6oQrxw
ZnyBZQ3/Bgm21XOF5xfjlI8F+YMX4jCiB7J89bF4bK+y7/vKvcAOSeI9d469KQxN
Hou4yDV81tYoDbknkhnOTPDCn+3rVOLk0wtIOy09Dq+HGMZrZRov3yRxDJUx00Tb
ToNsTcvVqAphzt/yTIzPtRN+hlspSGJMDRrzgyk7b5Tl3UOMe1wb/8yb1ZWSt+bn
ocsgheTtSD1U/AhD8B/evgj+/PPcbzrYsIbtDqLbi7W4tR384gWVjXiJoejpJew7
TVixZyCwImkKWprZewbVggwQ8gSyqx/5ed8eUBOvrXllp50UG6FWXlwA4c5dmLHk
43rv8oNtBtzKuAImaDIUQybugn11zo2woLZKSKsHBea/cUGJFnqiaxLHpTowhUC/
WJ32xnLeoVdXG667J5E6KttnHoA8a7pPI2ZKoC+hOMdHwilabMOffBuyNh/Vtxty
ndl0J4z4hXzRkP1FCaitVpQUT4Gqu9Juvn0PsOJ2/M/TOihsUSGBqhvnfwBFCULQ
mzo2g4o+GoAPydrJsz0KfiG9hAwtIJUYsH8c5WiNZ7pQr7AU79pEGt1IuRktA0/e
dXgkz5QKE4MKdPRqv84n+xGEhpmre/B9jIeNB5TvJrqbLEFEAbGVPl50qj++eYPJ
hyh0QqIPQHvcZSWIZrs/w6gbJzKkIKmlV9wd8ooXb2OnAybZOVpaQ5s2PXFX/C6l
GF3yxHglFHPli2T2HknznWWgkjVpCk92XHFjO1TEN+67ENxN9x5mUvZlnK85NyBr
J48T+lP//UbJgkQTacEql343cv6HVW5djz7nknapB0oMwdBWMo6o+fy419JaS1uQ
hKpVks3gmRHG+gsifT/c60vk0auMNsHc3xzYboC72rtxy3ucEdCzZSq5g6sA3KT4
3r0B8/BtK/ZFDWvKT3FQNSB8eavGsLlxLSr05KJZyiV7SnOXcQoFXdDhzQTSaJQk
h4ycgtR+2ROKi1CfBTLxhiyiiUA6ik8QwrkzeevW2p3EcOn4X2qB4JI8pVzjCQlI
rWdUrn1FwR8QZxe8cOSU7K9STD9u9MLO2bm4oBZUwEYRFXplu1efq2xkbqivDgw0
mwPOjwsyaVBA5/4V0XzMdGJ6F92LgYusOzaYa/jk81nJICYYnnJ26ceLly+vqfmN
XrVqHAhurdGk89Lc24x1U18DeRts5QOVxumBMrU3zpBJJwGr7druKXIzQee/IaVb
U3QGCJUkaVWSJq1Wnsrs/V9e2f4b94hAvcCD0K2h/4jpmB1W/KjE88+ItIu9e6MZ
sa1nMo2c5E3hzrOWzL6zGr16miFm/MY6uablrJxhX/t9L39xUZf8iGHYngk3qMZH
WoA8XBZpw7ovwyZY/eYJCLJqQBCtAJ69ohiCGTy+VRXXKzPB6MNzX+sSWmJe3wtL
VnEpRXs7Vv8eoVaNCKLGJw6Jp4T9S7HS0WKVAMtQbapcQIxPkqn69QxnSjfrWjh1
9OApO3EsM4VEU4B67bBruWdDpblijLRtw4xNt4zCHnA5UDFIREVHjsJZIlgK6tYx
ZgdoasloTuRryBdbKMqpg2bc1X7IHu79HsFvv8RgUIUplarJ0h3n2rYh9YCoUVh6
o/W3Bge7Ye32/rtRMDeqxdtKoFpQI2lAJGgFihUZH+7BHw9+iukU+JpsWAYrQ8Cu
PHCZmNII0ZRo+oOoKwavuj2p5xPPzcAui7AhPCiYemjo6nXl3dn88wwSMV9VpZsD
L6eHA40dYqnUPU049u6rP6vWK817vCzsXxYPV0tj/DuH+mbFFGwLXCN0rUoHs79P
j/m33ztzHdwVEaFeW5Cv0od0nB98jNW0BBlEZl0DgLBh/ymSnZBiMVJKBhhDvW/d
nR8lJA7MZQuR/zIjHLFCASAnPrfQU2wMEeJnUVyNoD7WOHLfSWr2WhBO9mVRp32+
ib2QFDLBaA5chmbDL1nlU1STOP9hkxXrg4uwi0685LHCMuDAslQMQGMiyl22/d9d
W/b+xRmk5idGBEeTLbKMevDcVnT9q/UsPXQ3hDq7QuEduIUa9NIOXub3LropkZh3
k9K2eBognpxlnZ0oJcfH77kXn0ihLK3Pxev+iJ6rv9KLWyS/mQv8WDe/fl1YKyID
LuQvVkGLKvkhybihdsA8tZ47mxhg51weXa7dMovjfXK9m9eVntM3OfKS1lW6z3B/
bpA0qCmDTjG6VskFNTEJ7pkLV/mYlBzjQw7jfsOjN0AEm45JnbfmNUD6YUR3Wg1x
kKKA3w+rUxIjY161BmJ3/J/JgPuqEzgkn5qmyMy6jguFc7OKl/3bkaTooa5GOEQ/
iH35/+nAe5RWhYL70SHlTSsS0HLRjCE1vPQqw/tt4hti2aNkv92QSiKJer7bFYWs
/JsCO67B5lREM27Y8quNlGoVba5zGTJsDUeQA1187lU5Y/jIIziZrVJwPBmI6NRx
6j06R94CFSRY5Sj3ac3onuEBSboWNsW+3IyP2Dxj8hQMtYZ7N7hQt64/0Kpxia8U
7nx+DhIV1fN6lA8jBe80NIXBpdH/EPTtqHrF22IXqgARhl8qcHq+lnImex1lCp+C
wCZdQlZYRYUfYJbd1tCZ+xvf1uW37MExWwy55Sc/3/53uXiiYd2OVVCEwqbUHnj8
AVanWEAKWC2hkHckYK5y3tew2uAfRdoUcWBrBTuQ8Dpm4ZIeyVkvQ/l5uWUVzDUt
19zeI72Gex0kM4u1HnuW+yHoYR0dqUgmyQXcU19b80L1hHzuIAI7e5vgiaWlBLum
QYLrT8aXBOl8Wer/obFnhPbGS1u/UhqK7t6jRPF7eX3J7r1VtqjtJR8fJnIxaRsb
zzGpQ9tt/r5+ghT8fff57A9gIwye3d+P6jXT0WAeQO1ckBjN05eocO0jyVuUh18G
hKH9xdlQIHaZ94xZRERNSeOHtkNVC2+rpal/oaOvTBXfiiqpXrmTL1G9wxtK4P5+
RqGgKFkiKBcLsDitwxLZ5RUTBcEV3i5zexbVrMwBOQl0xSKkUH28gx2z6kax43vd
Jww/5JI8ixpT1qRZzLuYr5Eee2o5UbdWKHnvhBBmPo9Pf3rWuhk2dJhbUWBussBE
4Tvmmy+Qc/itQUi/1WO0QdJzwK0KmeQBNrEEEgCHSofVUahG3jlPlB3NmxZSpRgT
PabY1gsvGsepmI8ibywBlu2aklDTBpbKpUoglQUUnUA8zqpEi3ri7pD1ZaOmUO/R
f8xS3O7lzqWmyPkkhqxXOjetJa9xKheqobXpQNDS1Xxehu8jztM0shjAitF4rdGT
nZEY0GBbcISjXiFPzBETuroIb+Bi6V/fWlzZakBWU81DNp1xSmlj4F0tD5VQitPF
sr9vwqKwAQ8lccJf4E3suI+EQEMKP5/m58i1FMo55Xkc4r4Ta2VhfB+r3gEmVs1q
jDy/+DqmGtC4hKwXVi/k6AcIUhVM6kL6ahlPgF2hd/dAsxopyK+9jfeIo5TyRyGD
uIzIMQJQXU5oYxmFCKHtUE5dBe37xSWHj7ICgO+8lKUT3txRgjIrwn5PdPTr/4h+
fP63UBlUPUNtsY57KmbdvcqKsrKZ1unPzITMTRm2K4aulstp9zJF44g6ZAczEjm4
mIBAyGul48tEWUVCtdBiXbmMUPDprxhl3epjgRxPD04iamMBZRcSV4Yozqn1G6pz
F70enr1mCSKmP0YpA+D5aKSiC3UPX9InW23GnBMFSI/pPpqqt49+fr+pF+uXSywa
TeeXc7IXuQKxXY0DbvbpLNxhu4gOaBep0aoeiSgjKDRo/WMbn4F8QnprMOq/KUF0
hdexXMZ/txlv845IhZpGh3X0G7TlYPWur9jVqE8fEjgBe66wwdRQjm2ZXObFpISo
xaM443sHZKJ/pBMVDgS5ByfPmQ1smgxqtToLC+I86qVWTvI4w5mwnapnzZ9stY9k
HAgnDuyfFcZywAqMjbq9qxqbcJONpOBxYnGgyQ0rS4AgZDObaWeeE9AzjtKdqFRP
NUgtfVN057og5J6dzlzMlhtDYYI2iSrHPuh0zkj6VcAGVIoTuWxrVuTMQBTViy1h
G0O3hlZTwa1o1xz6JKRIwGlLj46bh9UkJgC8nUrps+Fgl/XHk72TqeMY2liXYKZJ
gL8RK4G7cSUi+8xZS2tZZJh1AwMk1EkiuND4lhzhiAeN4x9wfbnjfxszQ09ob7eK
IBNN484V/bGe32gb0gEQ7S+fp/Sk0RiNN8OCps3bar1leYVaFI5DAywBLnrD555b
iEbqYxktIYKbDK3iZSzdBUQObiFZottVQ06LeJ/MAVOIoHms/5hEWPr+c4+6zUgb
ph7DJ58YKMFc0CFfulhamVssX2qQ/hdsfBBtGbnZxyiWBaU1yaQIRiUd4SQy+1Ol
xSpx2/07cKbORlBoazLidN5NxmmeQCpLY8UoYZOwoMFv47nUZbaFyt6oqZAxkygT
rTQaM8gPBmsv+4p7nIFV9Fkoik8Mf7Or8s8opfgO1YERuNmyXGiRurEuQHrSz4D3
765aHCDJEa7sNZAYlcSvh6Nj0W++JMMiXbrWZeBilqtGS0rZmS8KidxQP9OdG3ow
ijFi9LZR/jSlGlRW4nIdjhaTvvXTnEF9jTLQSqDkervsviKVVVSGbA9ZGjCfjCWU
N3UBySDZNyJWLPtLRLePIF68VFKP0w/rTZJmF3WurgkzitU7YOVS6Y18okOXE8/P
vs7ZpSVW0W7vZmghq22GIAFys9mLLDUX2PgKroAIs2gz1lIirfnOQ/40JaB6rEjq
ldd+/0qIcL+qtj0tolbigFDOOXelLlyn7jYdAn6jZRzwBoBkQkh89cmNJb6eImZ9
Lxl6jNS6cOseMI80faSQ3R1Yb2/WJ1due5Im5nQ6XzC4UhZ99YMN1qI3Q8xComAZ
9CYKtjIzEncJOpRPDObyxh/tsTSP0m44+a1qrnr4HI+KJnkloSH6HM00vncgRPMX
+i/Ycq3Aa7lZddjnRCrSdUDfFdJYUuafoXYCb4kF954XI76YA4qyyYf6+UFEoKQ7
59rvm+QNu1+7Qzmo5GgsQbccHgWBTHHumlNjyW/jyApkErVBQw80/4dnTULpfFrr
7rIauze6WbQQpcsrVWA+LUuP8fSe3qow/ZH6TxOvPVJNv0BMCeTz0nE0YuAQ8uFF
HXo4H+ENDi9bfPcIFGo12q36ca4FTtESEPsR9cYayOaXeYoWIcmUT2c0FlU9xstV
5O3IVdfQXAjdxN7pi7tPfXdhLbSb5y0DpmaqtAFFZbHMCbu24wXt9sGyj7vrQST3
A8qYwavVNfullRyU2uKWmjtIqru/ZWv08bbkrXeSq0gBNQbxH+wcRvCa6utb6qLC
VTn2vaBxVpsIcebmz3jcxF/lLRQIqZ6aqurAh78b9TJgjjKeF1XnkYZw5Y78Vxna
t/BovOG9iGYuY/aIK2lKSm1YnqpjTIsBz/cpu7pgnDrUuZqqAq0HUvomMLY5+YUy
mfc1ZXuUrLBU1ZBz5+AGLnWK1iy0AdrAjVURWAD+hoq6baGr9e28H/O7CxFilflv
0vXppCr+LfkjYiqJ+rG6RAf70NF8fdXyuSEwdzKGBq4WdCpuLYR/slZbY5eMujza
HhV1GZ1LBQko+YWhXRj1cbBbuU7KFRGd0s+FiKsnRdnkXQQkB+ZFUDkHQnKfq9JH
ucQ0l8Coi0+c1wpUbQIy5ZNvUJCZjY8Gauvn3m/zKJjFJOQc/ij4iN4a2ski0K/Z
RPpBEZjd5FL5QFVtYc3qBh29etWN79TPlxCnkTMR/e49op7574Z7jS6r6XY62nLh
qpeF3bndtCSgg+fSCXhRK+SgZf35u+MxuNhxOizm+CEx7mQXnNbcl+jDjcPhRPr/
RnSt24RT1HivwmtzLxkHb9kZKqEmdT/3kqq17V5CZtf6Hxadj5Eq651eDhxc0hov
NZt1ToV5PdZp4KTpl3qdCB5pdcbY1yOWqqL9DHAJ3yxZVDLFn2DmTP2mDqCqO1Ot
l08Z88gVgFrsmxWFMv1JvaKUB9BsALJQ60BgtKnwPsTn0sMZgNJR7Ii5nKkTCfWm
0nuEnO24vCdatfSycot6LKPyhbVmCZmyrU0TfMszeR/aLOZy2y6yr666Kz2+hnUn
tobPMqRv8raOZEC3g82IG60Z7ScyLoVq1ZJ5y37W3L7iYUFpi2Oiu1bM/r733lUP
afa4Mq2/E/t1ZlmaKT8IT2bnTapO5hjk3d/ooEx01z4zAAp/EmRbOhwGSfRCpkhX
A3RcuoCtmuG8WkgAGkxQ/RrFjMEXzOLt1gHuz1x4CrBnnec6Tdqmb8uM9yvxD/Ia
orh6DRwB+f1fTG5Ln6vRl0kpKLUVh9xOvgGtJfWU3nxobXfgFPbdJfWzj6UlOrQQ
IEoP5ZyH9uMX8a1pY6eGvfvzKkD8639BXIadL+CDL9FOPWAuaRgXx3oq4mdZs9oY
RovbuYlpscwNCRaoBfs5NTUecf3je3ASXe9+rpSOXlTqOBJn1IVThtPlPYH0sX9K
KDl32J+CHzdfqM/CuX8sETgSPh0oAYKambnK27Z6LAp9ioMPGTg1rIqvHt0sBuih
AqRiBB+R+gS0Km5qU6vRuXS30IedBq9SFf525C28toGqb/Ej9qsu/8GHPOvtSH6J
1N7/fLROinhbN1yZwmE39QBw0zYW4wg/XKIda/lI70Km8U5XSrqiUGe1BorQKMUw
y1brot1sNkgX84UhMP7iqisaEWEo0tcYMy80UvliUhD/rOyD7lN33zirvP7Jbzst
ATubueIiCeLHilVfzowJEjNyncB1qJGiOwQwdQ71ywi1dfsG/qvGMHRPc68tiZD7
xvVdHRPEJw7M8GtW8m3UUVIVsrs9P1I5xJbhNfkVQ7BxaX6ZlDZAwQrOsMhZf2pZ
5RCSKr9AiUv/R4bT44PB7Jukz1UtPWtTExa4aRrmBSmCypwMN+PrkbmdXIpOn9d/
Ra+e9JNMeCRDhGciI5bze8rENDlWKaHCLFb4H3BhmGVsAnjbwZHFiFhotB5a2YtE
D7WbkKRzzfjcdEahm164i3fsXlH4TTV7+Z/ld4SElP8Jgc4wCIaHMMrmTY9ly/Hq
3bd/4w6zklmIUnJjCtLjXHvb4XBFHwuywQfNd6MpnT/WYshM1IfriDDyaWV59sUT
I7TsBoe+wT8q5AN8m0mog1rpDzyeiz0jmoI8/YdDGIxGEOcf7UH8BTXC913zlVzt
lp2OdUwii84iiImzaHPZr/Pp6AhhGlrof1mdwYpecJsZujohRG8q0H2A5VUaoQaf
y+7ap4kIrnnQbDOiAr34m0oj3haz9YHoiqnWtP1eSJomwDsIY9bXKqqMbTRv4QUf
qLI2mljqiEl5FEq1NebI+R5ho9SI2LJlrWAqCGdhwVN92tOeMcajA/RokG6Nx3tE
msJJxE5h4RVpICSAzo/ZxKtBvAt3WVdIdp8hsyx3S6Q1SOzTGj7wbI3DzN5RfUkt
GR3D0WeSGtNm+nj5wA5FtVBl9wxGzsK6dNLFgiis/vj4+NXHjHKm6sk14FZTeJ/y
p3pImN4vDJQCJHs5ykQjXof23qBr06lozypUViOb4BNR2u35swAmnPtUf2ZnVu5Q
nMgpp21ss5R0/D6REPKKSA5ZNclnCvRSVoxgCIIBQ9aE9sdA5Kr4iCK8jOOZ2UO5
U+9W/IC5XCt+M2DZVXn5foEOb07gj8sffFFCbZljUP8cz46HDWwHg4pfXPyQmiLS
Md6Zmm5QcNZyapDBfEh8MG0IZicWohEcZWRD2myXS9Xf5yHN4X9bi+Qn2wmWNqG1
umrd+W966PkWwTqkD44kPwv6ur3fTlzLvf7Gr+5KDiAGQTjHaMcyR5lmfcLjKAbg
cSIXwZFqlQu1VGSfreb07kZ20CmN/Bf2zsqf0vY0rJMlnP3lLoivy2yaUZFCJRp/
3/R/wtZllAnCybpCsebjwx4TAdB6bRijJzxyh7tWhByvN1Qdg3+ma+qiwvrxeaGn
eJDbmAPGXZ1Z7SnBp7ronEnnB9CLZRP4PXmORhdMmwC0hzkGW7s9Xn1yXFL584SU
+SsXAiobdfCgAzo1YXGJbacbqAP6w+TNMTZQJ+W279h29xUg+HvJxfN7dwrxPpCy
Mr3iQj9rHskdEUjiU9VxsxZwoaOXiuXC3eX7MaQmKiZsydctKcdU7zzUcilQeXlx
rfYKCWGIqtxVock5gAigzSb3ie2aBMcyyEu6dmFNzv1oKUNGVt8ZQGmAvdbUptk3
ASnG3Cr8+uahOcXLAmHCya1wk6qOOGhcAYdLXDnSySF85vJnP6qvy2Fu8ElFrF8W
JLU6ZUpB2OYKSpXfvIb2AL01uqK3bJo5gXILUe7G/BN6wnpCU9ATjs6rySUhlPBB
esxehBgcpW20DXlhEmEt8Rr6COaRiNFxVY4jwBa1W7pb0KxAfDjI62sMm4uSEva9
vt0KUzkcwKAEMMEJl9rRpsmunZLN8GNPcSIN+La9kQR7AEomVbKqT+4Tchr5S8fm
ieMVOOHkEz6HYsPWw41YMraeuHlGZS4TY+oyQoTDmE/LWU9sTOKhGaEzYqh79ZPQ
dEIxbQzbyyH8pLk+VxW2dXaHdRPeZm7L2oVfdFucffjNEHMP/yqeyr5YlkAhM9zy
T3iwqDd5bsSPvCXsiaVEznN44KEZVA9sQ6HNzpXMdqyjAtJ/3IlgxoRRdJmSVIo0
nUMja2u2OSeZq9C82oOwR56xODTMamt2AlGBdeSJwAkudaTXGbhYFpakSE7NKNsS
YyzjNaLTFN6Fd4CVQSC0LYxeHzibVJiwr263982XFBt7cRN9g+KFUcByKgubPoPJ
POGX36MwNRSnbcb9yNrUGij84ye2O0Ng/fqRE1ydBdIJTtk18gxwSONUu41vl2BT
92ADhhgka8vIRDAEQMg+Q0l21WiqkSqiVVYMdaP/li7EgbKWet9SD3gJzQ8xWxBN
LaZaVFagGTcERfpqr6hsKcYawDgK+YJgGZvkaAEfcdx4SWZstfqDjvxUUJlzIWB6
mkpu63n9l2incPyqapI47qgl34ecIZF0jyTW3LN8M0CJpo/bVNJR+iwWABSe7+Tz
r47vLbmlcFknor0blPsjeALSRijUAh2zHqfuW0eVbyMZuMzlRebSAjvEVph7i99V
1H1rBooYbIs0H2py2nSBO9zkyo/TmBWjPT0K8eO+p8gIZNUh4JtBdirVamfzRm1B
oHay7JkKV12vXK79BYOnqU9ZDIbt5IgAmj2F7TL5Ejzv9R0rwldSszXWqwbBemr1
SEYu6ketzkn7e8d5F58/gQInwF0S/Kkkb0Uak7o5ouuIbiwZjH4k5h1IZLMnEbxS
SNm76XusH3UbPgOPkDjIW9ukIY5T4O0hXXIimhlNOEtVmO4WJM4DuexHMS6S7sXJ
P1iJ5ibwHhiFKhjIB4ThP2IlKO7l0ILxHI5jN5zE4uHy6eBcdbYhBFFvXENsJkRE
2Ck7rLG5oXSkEjRRokxeRt9Ek4IsSZENCJP8dnIk61KnjjZDBOyGe8CUAK2kgtYL
rzhNRG9bxcZqw1tBRlhYKgJdy8JgsLXFB+PIYgMOVkhQF6wOTwqVkZoKOVKO9L2x
eTemFUz0BDOMf574tYetBjyC2e7RIRy1xU3v/axtYQwE1jiJUvia2zsdtJXP52Vd
yTgoFnIEnN0xZNb5npzINIbK4vnbmCk07zUY2ju0fCcWo84tVPe28kYlKX9miIlZ
t8T8R31ohxOoAxey+9h0ThZoTvOK9WovQB42kbC2UWn80dFkkE8iR+efP/tPXTLS
FLekLE2HPh/k351BbBD1JGTFpY5abVgxqaz+wDRCtjmbEW0cQeW2DfrkdwV6in6f
iaYK6gjgbafbt2a2gwDVnXWN+bauNlsi8b4YD8ESSDNUhczUFElm6c+o7oxZRWZ0
z4NQ5zyI+8pHHJ+nV9kDsXljm4Ncjrsiei6RoAi0Ix0971ObaBWNDiGo6QGE4sjy
RGm69Cb26mZsrdYgt7LH/hVqqqUHO1X6w1octfApWotDCcmImJuLU42aupgaQsRp
k4tjXThbBO50lk9tomvUbwGYjc/T+0/J1OunKauVsg6HtXIuZKvgbq29t7Q+OJ91
f6TVBI2/mfRr9SExBDZvF+lsPV2hFiGwYrfE3ypo9NEMkbnw1+kEueMoo9bJ20dE
nOPx73QqkHkr7xX0czR/VegZAqE25ztU/7TXuCEjO2dV01u5eDb4XeG7UnoBU9HI
TYxFwmH2oiI2+8QC2rbZ83TPrOyqnlsXSXSYNerh5Dvc6xKbz4RuaM1ujBW8gJCi
sdAEWhzuCMkMCmyDLkTnSlpMvrLBm3/L1LT/mHI9im/+uFzozy4PV/P/cHU7hUzC
HADpp00EQhMkpp3PqaScxS4fh4f3wvKtJHLfwnHdPkeIEkyzjmdd4++kGxbAVPiE
0KeGpqUtkxXb8zvEst/AkDDDr8F5oqRHHQyqltPvAoiaCmQk4aWBvJkp1pBgAk8w
h/Asey/Er49N4cHaKL5hEWks3bujFu8DW4vPVh5ygE/dZ9BL3+ojO5RhmD2fITJH
yBog9oCVkZWBWJON3cv7oJ3aDJVkyPV8eDykPUtVLu9GocXVNvU5HBPkRtq6a/ff
aeLxSiYJr5NzG7qAY+o4DHR/ePIc6i2GESVj8FnoWLtdrEylZ3Vc7n/6n6M1Ulod
7uY0koXjOan8LQMs3sf63GQeJJKOOU0fRLneR5y1ERzgsDIpIuh8mKvAG80tMYXT
4Offm5BRF43tJNlRnv8H3GPp5DxehZaRMIZxB8yyNl3DcfLx3IQx9RsKsLBicE7A
gVjxl1pehpaqmRXtV0vYT2Hy6z44i3GPOlQmBVjEcJPQVWIUtA30yYJUf6v9Mq2N
cEwZHtjwKLIy/I2LscrOVh1mov7Zx7uTTAoZKjzBbFkkQQdbx9ROf6hW+Kjdbtam
gX83Ab2fCK8CGO34bBn4LomNOM9EtqipuNZLXbRqHyuZCi5HRqfvLxf5Up+vqF6b
nceVagv9jFUXuEQ1hughoqHnwtEVU+ag4wruyyf1bJqB2jjSGZnzl5u+/tD26fa5
QXyI7ye4foFRQMXmBg115YEG27T4KAfBj749Z7Qg58wl11P0M2cRAslViH5B2Rup
9IRugTzDMSnCdDuJlrngW7kM5Jn8IYtz+UajgLoUr/fsPWb1Pfi6hKfYJtur8JwS
R5A8D8R+VO75SJCscIdgF284SB8cEZfFPaKT9zG+br4gKJc6jjNeHTyeWzl/du9k
yb9SnfZpmYK1vcO/wilWvTlKuSp0Z4hs4Xt8FOxecAbyIGJUVBGOI/k5t7zNxtg0
FeZJ6X4MTnhQ3mgEp98848kno/WIqwJH0my2DxotX40AxV8VfWQioH9OUP2TDfwW
YO2W2+uWUVrV7PGzreSTVNb0L8I9V2Cp8PqFavUBZ4ZafVadkk+7RKJL8NgdeTJ5
D2EKLoQkMd1mqBoj6j+gkOpDKu1yishNpmvdffZbdZ+83ZNL6KdsN0NABWhAdMFE
dxqJWVAZZPAtiUAfiFx4C4vR0Qr8urmJoiQhxvqhhE7mtozjiGbikoEKsQNkhlk9
CLKnhxHiIWFGfDnhTgLVgo0l0hZqYA+I7+gm134dgDLis30Is/Mi5sf1dU9LRSQ0
xDE4NTs67XaWDZde8W/svB3Ot/tqXj2rwCel0vkRRN8LEhgxxJ7VaBjJWCaF1CKZ
u1AwwsIpNP4fPRazd3XtNpwYLNcXKSV3cJnQQQ4WfW2zO3Ga1v90s1siBwkCS7lU
5GvItg1k0TzyocH3sgJj+XR3br+IkMKjpMKZcdAA7gKRWMdyRxZBU6pqgDVUzy7m
WnjHn1nIexo4tZRv/W6BFRpKYETAs+b9qeGD3bEVj/ZBSs7m2QMCoinJ83T5X0wR
1mCvIKBVL5qesmQdn5ZFztTf0NiyYdfNggzHS2xyKt51IyQcftT04cFI7FAuPjry
NEr84bGvST/OQ5zFzje3Vfy1MfaTFxX447R9H+LwDN/q+q4YpIyr3iMpvskdHLT7
uRUegdHdxtDOJSz0OjZpKgFvTp8m4eqnTZTJ+dq/XUf8Wyh2sKJNWa4EFraX5K36
J6Vqon8P/o7uNQRgElypxClF9xvUC4XbyILY81ahehrNzwjHvPAasUPSrUKsBN7i
m7B27Xr4dAyXpa8fScpg+2RBZBhl1tCUuEAiX+wit6/VlBm4/JodlzUVYIGtvoND
p1A/v46sQZdImVzF3DbKSQ5qd0A7prlkW0IyixMZI606c1YiDIM2SnvA+ODTTaXB
wMWdh888zWEjmpW52/BPEDOj3s1hJ1JeB+8GMR8kef8kIuCKYKzrWemcf1EduW0c
rXv0F+LCyojx/ZQGVrAhE7KT7QproJ7kqJTU6ahOCFBydQKAwuZ69fK/490LNRor
+v6q+3l0Q36sE08S8wqlqDSl8r/zk7gkKddwcreYCXnYiOKB0kOam4KF4q1o023R
2QSXQxAbiLGuC5TSD2+ZiZrYboGvHNU/xQOllPCZL9eZK//5tf34jbcFaCLHMSMf
KAswGpD3XHuiiLdCA/Uwc9nQ9y2iqwv+ydN5i22EJadd0mpgtsyjvBaEU2Okj8Hn
NcRV1AovvELQ2cDueJr14vZ5jBrsP8TwBkXLQgUn/Z45KawwlHvhqttjMeCNr7FV
MHMRQB71jd3NBUBwWEYGkzp80tnYimkooDpELSG9cbyti6RVrrvQBiNp24vGoykt
feakIYQZGIUI84kkhBrMnjF7IZ4lE+VaId6h1xd4j5c/l6olb4lKB/hDsEFHJq1C
MKs9EeRF2pIhXgRvoBnhLGrP+hhJwHjjKdTCcPeXUplcK0TNkUOLktEW7+tDguvl
fApuT3NR6pBPlHU3xO1VvQtLalkXzd0JwnFgsTjqF/46N6atTWjuT74IdjCVLQ9s
hF21RucyG+INAnI1FI5jQ6q/Xz8yXNuUafJSwSh/aY5caNRw73vYnh/R/QKgRRQ3
QDOoNuQZcNla7vw6ZKLbvk4iyp+XVUpFPpY+Xl7hCUKySYDw1FaOmbxssDsQQQg3
ZxxHhwAtBaoDxqvlsD8V37qQjXo1PXWLOJ+lZO0Jy/+sI8cu/9mEvVgNzuE5FvoX
ank2UuUkxU6dh/EHhzxyvKn3zw6ua2xS/VTUeo2Im5/71iIWOsvalgQbcMcEgJHz
FnxxE9NXGUaJ3GBiYxIsVE6OhnJUGp9jNu2UPDSetxq1nTqT4F5w+gECm6pCebO9
ErsYB9g3a9CD/96lURkwm6t5KZ53TF2Vw7UN2RYApxOsxBpZtHfb36sJBpjZLKJX
mH0buV8qkJIWGLq2eFbyS1TD4QaMAUacSOP+iam9V2z7fs+JffsrpDevKJQIh/Ms
2KNUW9zXueFALKStt9ANN30XlQwKtu0Bq/ZWsk7MKLJbeVFtOcBi9jmowbEj4hTj
UnQ32ag7pbV4zspxu3mOp51ZwAbuz+n8bjVo887lz3cQ9jLafyMPqIVzHBnM1Phg
SbU7WZEYTGFpcc4+674yJT0Pmfu22AvJgrldw9PR6Loe/qFZ6Ulwrwvs7RSGieTT
F+LsAZurnakXs1YGXhi9HcRy7kR4dEnI2ZhPpt4W8zWquDOHXQtpKC2kCStB4VRH
T1kEDiiQZ50G35K+TOqqh60s8AzEpBhRDrYeVEcLcSG6aA7s68NTuwP3s7Iv6ss0
YGebR8buCTK3vgUbbJXR5760Ij+EVYg+RUM05xQl+yaPghzIUFiGjuTCOef4xcef
oszVhIiDOdoSMp+adOIBOeqfsuowQEjuu0MBaTxD/wSzQ8/nlhC8yhpKzC7NfO16
udQR49D+Tp9l95DisGwGCnGoXaJKcll21Usnvr1AJ7CRfwNc96e84bIMl+8tdzks
XTAGgKhP8KcreWpNLpETquWGXZYlSCcQhLAKDCaDLDGivaJhc3NIeLhX9Wa99dPR
4p/pTAd50xghXS2Me+aqBp565yS/Zxq0BNbuwXBNRqf1CxNtOzUCdDnAJwK9904N
QQchnsnJ0n3RbpDGS7ro+7cJpqHPzQMV94DSWe1BEjsFzPnDO4x2iQjVMjHP4r+b
I+4ypLCE9hqnEJnlfuFYO3YBqXMPc6XeFYFh+nKa9k4XI4r1yPXc+bQvykLc9xyU
NslZ9pdxRTmAGFUJxxIkTFY9ALvGRgFM4qMT0Ei4S4B9y0NkKFRRdazeb25E6y2X
/Kg6V7xABwTdtUniZXOLLGu8fu/NOWObT+Vk+BL0XD+oZNi0VkJFphtHoLa/oX10
mH9qRG4tgrF8ars7Z4KbcsC9ScIHRNbrbWI+BuLFDInXx2kTilI2gqyiKBItqGs6
j2i3VKSDHUTmrg+O0gM2LdVPRTDUGdSRKCmZFBhe04WAlt1Ow0XJ/J6NYUsEXsZI
7uM/pewRF8GF6cyh75cNWTPC7nEzomLK4xuTeI3e2sVoJNxDp6wYvXk44SLzXVHq
c0FRs0An9icnS4c3VCIuAzhCiuRWsof63Z+7z54566dmfuEjR4cwwibhY4l1FZBt
VNGluGi7OqKQSEpznCbE7utagXJtqbc7W1+1rWqhCF0rCjSSR/2I9Z/Jac/LyS/f
BZGHDk4gkp+qLhPifwgmUcPskhHyglYzSOyJxWnJ9Bfg7XpRm7w8VSeZEpFkEcaF
QWhbFbZ6xguLIxZMaMNLGUQZlEhbA/x1PEB3rILolJ2mQbRX8U3+m0mhU6KQq0dG
FMJ0hWuRCkPPLkZ8M13T9QOQ1QuF/LWO+Ss7sBDtoTvANt6egKoNj35HkkuPOt14
XVBkqCb32xVgf84DaQiYMFop8sdClMBDwgnwCv4dNTvCA7SC8k8YLYz8Pia6v47+
affp5L00C91D86uH8CL2iHdhojeqe8SJvOxqDIntqrxQxeZcd9nv7TGfzrZjFvaI
E1jkMSqKhrIFyUMCvV82t46xs83w5liEr+W1SM/1C+ng4js039whfQAerLXd/Tpc
xf+X35qqXipIx1BNTLgkBLaZygP1H4fwxq+1WnRdrQNQF6sR9emPInbvEABLjoQL
49sIa5s9OKEfQDUwXxO3V3YeoCvrJmSWFlBWDxISbx45YOKDD1uT6Xhyw0eedBrr
wHPZRsC8OSDbdej/ygPiwPJ0JBun/arZ3/LWx6Z7POFkSZw/rUMwSQQrjbhYFgnJ
Zp9hcWlg6pr38g0CEBjUewkLwOhFFOig8Dao2Sw5HpVBpdglI6AeG5A5fkQa9AxN
2P49zA+FxOX6Aq/NJTzMmIFP5sNvAD6W2X6yooSxnFyq0cAQVltDjI9VzcWSkyoZ
gNtb9iMgif89pv8uMixZYIZhXyrjPLEcxDF/aDViDTqtrLC3rJ+l/aIkSGPCe7nZ
TySsyhnXLGlAXNTkejYeJROZp15Of5DifwenEwvxccHM2drsTtcp/1fLpkML8tAZ
PuUamX6R8Z2m7HRqvRx3KOTiwQdcIaeUhAngIE2sN+uxCG7jf3vlTn1P5Xl8cfpP
w2DiMDrAx2cKkS4Ex+NWAKlkPxqfRqLgAXh2LMMaQgPzuQNFx4XOBmp3kvnKndpW
hP20cmcYGIy04/3fulPLrYmfX9SxBnmj7bHe9obHr6Ypk285QanmAqt/YGtxlb8i
2uE+go0wM94Tcy8Th5pnJbQHWvUtDTV8LLAPibSDM2Gxnv9DRPmWoJ2BLKY6haVJ
TLsd3G3xCXFYfIyZw3hIVZqnaJAUKQNk2prcSIxK3xnRjXpElj4pWcfOhEvnNk4P
IYSis559GpgX9BlcZBcL/uZeaUZrSXHw5Nl69o90qXRacb+nXtZzXoZalRlW2uyf
WFpDth79bGF7J29lVYaO7QMeUvABJPEQhR01V82pwN27HjMb/apvjtrrMCmq+QHZ
RFakXoV8lf94UalSNvTCWHRSENCHL9GWxGD0U4R7VxB02wzm4xmffLhfYiowQil7
FpdBQgFKOaqvdonrVXTm2q7WaPQihtiNdff8dqAHmIQrvjVhKGA6jymt7SpZb2lD
cmg2+0m9klFaAYqKi94Zct9o7vMDbTQJcFTczLKdSkmocPc2bZwWBJfzKLOqB98G
k2fJe2/76vBTQmFGjy/MphMTXcFb7fd3gli7RDT5WiM8CO5C1E13yhMWJz+LI0/H
JBrIy6X9xZ61NNFBzN9iVC6wuFoj03G6bq4N4TTTS9cMDjKa9jHg6yhPVCt++Qe8
WwvVf+7FHH7tu1gVFlWK5rYipP9kn/7SrWw3Uo8yJRZu0qVzOBD0p+UmvE96dHzV
+bKNh14SYkQXaFS3GJpiJH3VtcHFDv5N9r0+a5hh+P1aM3CqU9FKgfiuR4ty4Gh5
NmChojyEf02UDkHDGm6CNp8gZqqv4HPJ26bHpK9CkC3L0a5PE2/o+XRp8zHiYRST
gglLWFMX9t+1B1aCL2Ss7grl2pofhrwqe921rhwi9GIftaP9gZVByz5oH9ZUQQE+
Z+FKLcVvZL8MuFMd2aAyJSXbYUkkjT6Wr6ZCz6jEASpBxZ4Vh4n+mTkWpN5n02zO
nqd+u/0m64uNdQMxz7z8jL1GsYjFZi00HZZNXF05fUVz0IyM/FClltblNub4MKPP
uXFahpLXcltJ6QABgUyBqNmdueCT5YjaGnHoQGjbIfsQHvXrDDX7u2qlRQ/KYMm/
eJ38nQWd2DOSsIneLipnTizwyohCAUOecABOYFpEbFvJ7asdjssYERwq+aORk3+E
90Ips5McBc9OtCgUmp2lXZiiHq5sFu76RRS/C1tcrlPzT7ZeMiJGG2QmrZXMrCSB
sR6yORPWx4PRLFQ3yvZ3F29wak1QJ0+qleyK5LKfhtGZELIo27ZnNgigzhwPRaeG
0WDwZ9Ta3nTG/M2TCM6c4as2aBX7BUUbfSJdwavaEFbvFdugPPlvTym+ETDT+DJE
i71+qgC5/ySjt+/gRd9ez0yjlqnKrMcV+jr75PZQOidcbY6xKk6ArkYgo6Xj4shs
ML//Y1zZx+Ort/vmLIUqND7g+loWw5gOk3D5luYvw6YaG3VuybbWWFNwIWsKqRAk
A35H7dcvK7+l7RfCl9kIpU4s1abTUCXyfhqFMF0hEE4xz6mVZ/3U+pCU1DDlzpdJ
9Brstpih7quu3jxAIQ2Yu0xmmnYS4T0hIRC1Kv2v6DvIvzlBDe2tevn3ijCMGiGs
tMwRAR2/pk5DtoV7DElnusOwS/OuCDGJ7KzjL6rgbhGL8x8XL4ngGbc+GbRnGXxG
t4UfiKpG3NCM2DKjCtW0RbkHOCuRIlck+Y+y0NzzRr2XnbjFxyqdfVU2yUMaA+fZ
/NlvzXA9ksCR7vNUzQU2y+zDqZdy8uIMH5dnjbfxPCuTf5O1vE+FcDkPE6DmPj+0
0go9bKbtq1b7sBb2f4llukXTehmm3/8g/MLKcwsKJAlLL4TUJcMMSVHQRvvKO35O
7tvD0f4eMOKKWoVdhU4bFwIBZWqTXCycBHoYqfWVgXrfUBCpvA1qnCp/hoH0doPa
ZtpmAepSZ3A3Vui52i9LG1hcSEV72P1xk/ify4W/y3WvXWaXFd8BOCxCZ+Mvj/1c
fBjDo/Vii3e0jLjwzCh3VH3SKlRnco8i6yLjTQxbU1qtDHA7rj7jrjAGgXOjXNt9
jtsBfEAW40QuzYfMdTtH28jDscCawXVRCN2h5wgMBgANukS8z+yXguWdXONf8FF5
4R7bUec11jAQTXWEB8dX/ZMQ4Swmlwl/HHKFBO8pSOhLUDwqrAOKxTGqqbxmWBxU
ZLy4INyYlceEI9SNHqQddwOQuaUEcGuSOTw7NNACkaRCKZopaPH/o23ZdNTDtmuj
G/rMcrCVErAMHfK/nFfdlltuVQg8FSCY77MzIhFiw6THa/GDnD/qEPZJ6SrK6Xj6
yrWc7LmswaiZ5WCRYPV/XTRYUz1mG+gznG9K22FgqmME+s34BkHud/tUDpliTk8R
87ZVZcqyrVqvh/M23mWR2HxP8RhtOlQkmRBqgbl44JwnQjiBva/CwNgWj4+zls+S
t48XIc+1Cklkd8a/7JDbVtkk+q2L8EngIGGHZ3deZEq4jHD2syks4Xzuur5yuyTk
8GG1hdENmxpj8qGXRU+2UKHAQBQtwkoGL2SG9ZwfPPMo+Fdg/whxoGaPbIFtAPPk
U2l4NHzyxfw6NDowCROeVsgvS92LN/OkM/woqzglfDBmXfRLE5ul4qgbHRuqTQzV
4k1u95urpd5UP6hpZAYriFE+WnR5IHXhulDw5ZPqyK2PObdUEc1dpQrwyHav0TJY
xfgFC7jJy6ZTGMjSy8LM/SXqv8hoXQ7aMe0rerCS22JeODxBbaLFiPFBhIebkvQy
LcJ12XW4NHfyowraxjnxH+sSkSO8FeQL8SZOXMlB+rjWSeIiGPXerJld2HlJrYCF
hvfdSu0Br0ltIiAcuUnQLil1YkM5pRKiDwc4SiWnZnrXJCsBjrCfK8y97sQjQaSn
8UWkLB+x1+UoV60X3ve5Sez4iXrGTacNN4EARdAzJ/dmE2qtXsYXjlc/Da4ShjW5
4ZNwmuFgmT2VigEeB4PZ2dsO7SR2e31SdGAVtCFH2qI7KM3O76xX8QBZeepxEng3
4tmPMVZ7NGGNBe1TrZKYl9dq4w3r5JO4hSrliC4T2Nr3+i3GG3k6qJsoiQ4ifmI6
XlFHUDApZkvK1O/y/KTxZFfg1T0k9hdPCwl1ShVZTmn1TFtmtIzvFJXU0mE3NL0b
CwUbS3WhVPIKNS1BY9Gz3Y6mFW2lhxLaUInfJzn8/9fyZhSvwOJKz127i/cv4/ZW
2ETtLuTWO4+bluYv86yPy3tiAI4IyJ/jupJ3TOa2THC5afHbFKcAqAQbXMzCyx7Z
sTFYdJW26f2EUTPyol8slCUhgbpmByjMfdL7oRZOIGm66Qs8EvEd6Ya1Mg3/59Pt
idNEZo/XF5y6bUnkBcpUqyJMR7BNBDEO0tcG/0ZhYePWXuJfchfAMkrPlUmCHmOw
bm+9gPEmuglrB8g6vFK9Dcch9QJQJiJV9bfwaO8yDiw+OavmlU9coJrhdIvEsF+L
yeagoAAWKDUfmlu2syCDx1IgayIUhQzLydMAuGZbJDDMeqVs57zAxcJuUIyNHrQw
03/V7x1zCgxi+5Xyfvy6u5T/DtWCxOOt3SEiM7/E9UAHPiNMyMnCEv5dusi/9nv6
WaGInfufqiiMZAmbWcgGmiysuUAaeRWjpGK2K+0Msf+Vw7twkvoH7Lh+Tx7KAKNg
0H8B5j22hVPK5svmgdHjLofBSTG+O4mzL9qrdOMhqmtWIHDutm5umyWMhMRx8n8W
ZzcI9DyrcNeH/3awNYYAmW/Z0trlcRbKON3FiI0oNSKz8xGTtP14Zprx97ohL6pt
8/rqn1IhIMm83LWMob3p05oA3x0nMeJKLdwllrzTpdkKfkhidOPNFiIsBqtDfJYe
cSV8+peS0Q7WLkrieprGc3CHwNoceaq9LDKis3iFOyjj94ZEB/8UTf+2PEXuQ13V
zb/6kNeuDekwRVijO/DBWVOPVMyqVxRvbWZflpzYtIXE8D3Sk/4fSKU9vx9z+uU6
Sl9uZasR3wo/eJ0Jdgc2Uv7Ip8H3STiEDi9ESc45Ced4Z75UX9JEK/+2IdAsLc5J
WAe7qYc5uiuSmIl7XKafO7kZTU+dctKpl0E4Zbuem/iXsGUzhJDz++E9tgFTvKzN
qNtOUisn9173HTTL3eeepKflHwmcmR2zd7y6sLSAbv+DdnjbK1a9heNApPaJSoFj
0yScxzdS6C5qFTHukIaEX+4GnbeG8T49uDGxb4Ap/hN8Eekzpq15InHC5fG86Z/X
v77VHe5zN/ScT2CUOGETCdcBx5K9Pf+REWSXzcgsa/yhHeKyxu8AKfzJz8KOM1JN
O8Aah19wh/fwxn9mNRBFtfsSslmgb38QKuukJeMifT6WlUF/MS4mBXtsfNVWrrsd
F7kpMTFYXf6Q3bVdP+RWJQTVzcEJcVduhULb6jOkRD9QQ6ySsI4S681IwL821Acp
GVnI4rSnu5MZm2SnNxG0t0Kj50VpsgTJw+oBfJMczsrhLn+RsxqhdMzJxQgQoKbo
E+VljQzgH8ZeYIRQnYD6EflcaeI5Xpt3nPwBROVGmjnlC54g9aLYOhns+/PjOPHM
wczyNj4CaOcoSxhcFsnjENCLlOmktIK4SxPVOD8BO2rDKNKdGKkWvOQ4Yc88oGS+
wiM6EtEkE9dsmMRGb38GSRPo4oXQmkeIs2vsy5r8D3bS/or+ZMs3iJdZ6oSRaNQG
Uxhd2e6y9m6B4VOhdkp3FtZLdsatni1oKnmp0e64tQ8WRC77+DIRlJDN2d3nbrSN
/L59lUB6Xk57H099VZkJOPpktz8rWA3hDOXGjp+gdOJllusGd+Fu8chzrbHYDNDT
gU9Q753KoudNBlBteW2cuIEg1+wB2VoRLJxG4tF+5ql3+nSECnzGA0UeDpyw7OMH
X6mkvtqrnK5ABqLrz4YGXEXebjd2yAI+acSn/J5G82ool8hXWey7G5fAhotcjL76
7nNsfgDmfz7Ey3LqP9NTpAJRxJns2alFN1GBAl3DHci2Z4xNDotSWT5amypPRjXs
huUtMMHNdWeRajXw0jb1+mdwXMb3yeT3/NB19DYvn8aYGkadfgimXYBkavy6PTiI
nLQk//k5AZzyKOpqWUUC5SNNUg1JP7RVMLM54hC5eie6XrPJuTrL4EIdffLR5o3G
4YUy75F1o/DjVdO5SuFA/6FjZ4xFKkOMr6P8SbkvL7yNpgDBaJv5zrfl+koZuI0t
ROm47dXxeXA2rqmcPpEkolpGBmbnrNkdcOh7W5SZzt2Xcqr9Eo/s00HwrJ8oYDSU
mGQXoJSfTY5+J1GpIZjKXVZg5Xl7u4SjVtO4+ZbdJOoNmJEu8Gk2oXNRtsRuoEUT
P6iCp/b6QpMHCxs1rZ4vlDGwc3hFdND9tpE90xTbp7Xn/iihPSzXAFybrgTHsWRd
25f/xeo6JCuRNFVJt3uXYiX+EW0tElESaQJRh4eYk8zd6rx89kld93uT+9h5hGsk
NxydJxe4AnA742zp0s7Mf6MCBoWLWwuVajea75ONbzJaskX2OXdk2sG9GTjPdg6e
34tQdS3Tk5tpaNuzYLiRnknQNfNawFpbf56B0LQm72mV/L2FhntURluqx6QU8AVU
AJFTG0hxBwT0TJMizH4DaekCLEp8IUTPxfD8MtSSr+xAVPsFZDeTASR8vXPLIb8p
3fvy8ddYs0flqqKN5zTp3lxV5mZVOE4Jzuv+GWB3D5opRVNoFT/ZTlYig9zfCWjO
8fCwixfSB5omGg3JfQCwhvpmsc35Fa8wXf/yMKc7czafJyKCNwwTTSf0FaoGxKV2
Z5Hh12DstuZvDAqFdnwbRvsqZU4TMZQiEOMen7GWA9oSWdbsKilOzvfuhwDRgtvO
bJdcjrkE7TiRtslCtZyoqHvaxpr/8YTZHQE60+ruEDsVDhFLkK8yAxWcFvCabm/F
KSvtKHIUmT+hmGpiOhQWspNa17k3aTXXc7ycPJBXF1Mvgm1ZTCaZjT5AD65QOSp0
9uUubTUSjtbIV+NaMpApQEBE8BHELa6hRyGb5jzRletJBYyDjAIhT+zVCREmTNni
9BcqTou5k68XqoAQ3ugTw/2Xu5cHfOIPAal0GbwKk1pXpt5c9/VdANcBOvP4BzUK
2IU7UnG+b2ruOxrXulCQPnI8nCfKYlWABCuS8q9Iexzc0S9au4uShY/ZBy9WoseW
6CQgG4CM3R1RS83rF3Sa6NY5qFsO4BkfdBcrzbViqwIdOSucpswuEVUlYdp7rp9W
pqDk8UsGXUodwYVlHrQ9tBhSprdbVp7+aJqyrzzH3qMx2KQW2eHHgAtIzLzuPJMd
jyzFHMUvcZivBzWMiJ7R+es48+5/p+e516aCEv1h3rCfWSUnzCOf6UvsWUGJ05dG
MHAAf0uWno+Zz+xPuW8mlrvo6inFikgx5iaKM/05MhGNwYNyDQfCjwsnVZbRWZKd
mAenxvCMTIbBVB1Fwg05mu0qVztHI/4L/1RxwLJ6OtZcjoaPo33K9NqOiES6j0FS
dUB2DMjIFuMAC1o9biVQ+2XjeMNKsJmOCozOGUCNW3TQ4ds6XcLMAk3qm5F+g0/S
8hb6of5czWM6lwcTuvKkjQFOhuEde1cyPw/Dth+14dJ36NFhoifmJT0KFZYsbVPi
q2E4Oo/UogkTbjWfrGDh1ST4pxpv/Y5ZX7fglz94vb38Ahrlh/YHC5w5TfJg/pBr
56d/akVBFzbN/fQWJGpjH1QcooCmFFDbG1i0S56K8fKaSXl3y5i+W8TKKqOt3NAB
Z9gHLAv8yv0A2RDhrIaNt9aeHPnJ3+32+xJ/bQ+bKhDdnKSJ40pdz97aV6twzto+
601XWpFmtoa7KhFBQqqikLfsARdzWhJ2yKcQc4BFC4FkAyuEohQgqtVpTe62D5Mk
b6j5ZDkGAS4H337+PnUgL5Jw98HNXuTdY9Y2En1zAN4MPEIr2LAR8Ao8X+7wI7nm
wT4dq7/yb4UvtjbeEQ/UvTegK497Q/nxRbnvnN0u9axNc++DdmFaYBoiA3t5aymu
DOnkAQlYIrP0bNlFLxrCoc3iyJBHrOIcqgQULggD3YzsDyMOMUAzZiZD7ubphzVl
TUMMeEdhc3vDztNYjVV3gBPtO46OPTvSTIxRvGZ4hllxd0PkL7hTJXQBwd2lfaZi
IHVIZfkdcq0A4pO1CAKOLD9ZPY+DHIkM2f7NOwK1hhzcgKCisqYIcpgFwAcln0t7
aIWBnZlyhQbvZEAhkpV1GwVH7uAYeICSDBdqtNFndQtS5rhO7dJltXpyMBP80J0n
vqA46ItKnTdx/3LRPUK9+IYQjXV0D4WDVkrh+jvI0iHawWzpj5Pc+LzNAvEDoHMI
Dlh5FeuYeSqpNEEZpyrAQZ4Wn9Jjn5b7CyQ8fk0lTPZKICZmA8iCVGe25DUQC/Ko
1aUyQY46BrcY9U0kntkffXJV7yrg6UyimnaKkOSJLDl0LsLZYdz5qSR1+KgvUQSn
VpO2Z0iFFzx5IHpREvOjyeN9IN61BJap/GuUZKH1JlWUEHoqHCdiAuMzVYnvkHrL
jvG8tdS/7+ur6UMUIMHPlya5oK4+NlmuZxLvXMFwhO/V0sdQ4sOzDWak+W9mEvOs
ujsEdKfwJBpzGg98mOsJOlmMlsHmQ5sauG0FlkV8v6StpZEyfh/76l56/7rDSrE0
MWOUQn2V1ngMjIjsqJVbmeDZ+sq78TRKbfdgZ/zKJjjtC+NMEKQ3KIR5tzollGnY
v7Ov8D3jbTaCnM8zDzOawfOgPoO4cCHmXtc5cXDw5UurShIelio5lRSKpcjo3Lch
XSVvf86ASUQJvcDjGQRGiU9I7ZlaEQisEtLnXdZOPnndJS4p+XoiFzT6BXv3VRC0
h59ykAibD43pkKnpiTLIw8M4K4uy32uK4ldDK2L4u05Em6yu68k2ypqT3dlzD0lr
4x5GJlb9Poe2xtIUiHA1i8OG41uOuVcMfYqOwwIFnS3kliA4wY4qAKyaHO7e1ist
53v4UB/vBwV8LJ+xhmefMDa+d32X6yhZeLIGp9gi/U/k4Kmq8SdqYU4Sy3lDBQLV
mMlafSKvEkmlaRYukWQML3U8VDnI21IIoEZLZ0dZLAqk551S+ZExqzW1BspovFaG
gLi3lq7Rfnlr/YaNoafcmWoSoBf9YcdfW36G6x5RcAXzCavrmjpmvNZrB67ntS+H
bTJ2HKuHOS1Mv9QxWJfON/eNHB0VGTfP089H9ntgGVN4cdAOmGhurB2vQRb6Cs2K
AkbBxs9ccPN61Ncs+LAU2/sxILpc0gkyQ40tA95NnFFn2Avy7s61GeoBC+O8V331
hgc8Dh7ZR1ZTgrY1e7gk/1grn+6cY9QghU53y5TiTn0u+f+60ezPCXcJNZplMbMG
vKrugQggayc+cb9jAs90Ymm+AprqnooE57QaOnaKjQyGv2DJTQvyxBD7KTyzSSxV
HqyXViurul+VD3f2CWr1R1CHn0HYXjv3S5eB3LkwVLCAWslpwX9nqmhOgku+0bd4
G/WCQjgSjihbFR6//t/sdYua+HTsCFEOcNcqXAOW/K6ZNRJCCSYm5WbM3yxN9LYe
K9kaSl38lAQF95Xu4jdAe2FqX1HNbBqkg867Cjb7QtgRka5rbFy3lqpD5d7YxMrM
BxL6eAWPNDdF5l7CwAOU+8+O8DJnImoY0vq8CrYVPdTzWcCIYWUOsXUzk9HTuANx
NhDHqJUsLueHAlGQkWp3LuxtQOi9RUm7fyw0D3o1UGCWRy++MG76vE6Yf/Tk2NP9
ZaP1Gbu5Qi8CsdD8df7uFLKVyoQsXLnFJK9SRrGxs9W144+wL6ErEAfwghJkJTNO
0aq67pobx8OG4UTNM7sQxHNjyN8PRlObY8FWwoMzjNPGJSI0XXDG8O1TwQ7ZYRzu
dzoHs8cvt2Jj84iZyKd3/Fs3MS/NOFKhvGuRuv4Fyf1N6QyUscZMBpULkqvq23If
Q4Nd9ClA+VvZNAcGHuAxFyr6kbnCq3R1ISgkf+uW8jISrhppliIuKTUY14Ilahov
B95UaQVLbsjz6pRDjjzcKZsTqyovzF3mzWC5//yxoEz7Q4UHJ2obGA/lHyr5aTkW
di1nlY5+EzvmsQCNly7uW3E61y503tszEmcoRq3KBMglkkgJl2xB4hLdw2v8ickd
bwiJ5Ll0H4x2OY+Wg29KPYQW5ImjBdq1FqqMWJ+8q41209rzFXMACfDivh5e/SHe
CdU6wUtuiSvISluLc6qdphJOLzWiJwfWeEY4iR4/RfpDc97TJKjUaqst6xJQ73dd
q6AzCynaYL+s+bADV8C769x8o68Z/DzlejMBhCd+vU3BtOB1u8R+1M95kIQwYwbN
6cf6VpU1wkku+8dOUL7/JXtTohwyZiKQCPPQqtk2KafNeL3vsnjzj3fQ7kfldPWM
2VcwzpppCIxZI1Y4evRIBO3QqEmHkjE/6YW/gQlvH2bY6gs6qop6KDvII9EKOSTm
TpdgEsEhoh/azB/+QwZ1+cNRGlNXMwWQvNR94hBkGTNMLkWXjF9JQNb8heFyJ5iw
ks+yLcMgyw8SsZ7y5LX/JTxA4k3l3CQv/gDYVryteHJ3tkTJCelRHQo7bgVmxXu8
PECpEevvULFSYb8zOZ4zxPAVPkAR4XZ6FJbbsPzCmJuS420mL8Fs6L1kavnBUc3c
lKCF0mvbxMZAM143bVXjFKx9OhDeRajD0O/R8An1VMUcXWuYqJq7Hodz1OHFOsBN
6dA9eTn12cXgrQa222+XOR6j/TV/W9V9tCVoLBcDlJCTi+OBai+04QpHvyLZE6yq
WmPhDZjegrwjg4M/a+n3O0ynQzOUDB4RpyQtVCBC/ItVLSfdE+SGhKxjJZnHN+i3
4f2HPVcHwbWMaNSmIR1zHZEUgRARdsim3RwyuR/4ITMO3GrbiUzHUzY4wgruXMza
R7Duo3chp4udcM1UDimzxDYQKWOHktJ/pdn3T6UkZ/76uranRHbsWFAXM6fJK8mA
oNFJjWM2OkX9QTKf9DoRXe8uvJaQAB3T6J6Hgkn/fZJaFNYCaAYYdFKdHerm4jwh
A1pAkh1G8vwkAUBPmo9pJi/F1KLwmq1zAtQotI6IHK/UxB1kWl35TELSnX1ERTEB
0BZUXgCmhM/3kucXyug+XOz17DG1HebxoaZbaqy0ZXksGgBmdhEs71+IPlZaR1ji
n84jRNcWAoRQgBpv0/KDQxoVVrmIbR/EFwETrNOHi1fq65cZS2EktrnFaNx8SXRM
IwUFfLEjUwu8olkGOKeFNFoHH1voYMZuTEO9HWPMvbuQdUUiRBqwkfThsQRnUw9U
6+D4TFnL593pfuCGbCawMXWhGN600oSC2p9fX0v9eiUrBJe73C5F4p9SBZwOsWnB
kw6IJmmuhmQL/VSS6gvWCjg5z5wUmXoJkQdQL9BjjEpar1RfYcoI21Y3Q7Z0FUL5
W1e5ZiwO1L+xF5gAVGEcQeI2O4032MIQB9nOP7TxNXDFPTd9X/7zBzdo6j+/qKbw
xSjcvsAf4JuBVU8XOjW4ZtwjHw4+gXb4lN7hbyWbhdRfEtWxEaVqUxn2cr2HK9uE
idxODmlYbqEXoVkONAPDchkXQtLkh+iAz0uL+fyQ3cxpIopYCwDCFI9fZtM56xRm
TlG+sqCmiZZP6XACSuMInUHL6UW7GOPcSg5PkowMWvowYdlVLBR5pj7b+8l/F+Ie
FuP4ptl9K2UYbBs6SmyPBFK5NkombfayE0UyiO/PihQzwRlzia00q/1brEEO91Bu
qGjkA4zvTVTxtXbP1/CkBzkxWvgC2N+NfKxydXmP1SwbZDaSoBc1QK0k2t4anWg8
Wx1hoGE0FcOpxeLmoQdZGW9ySVJ1dAAOQs1bVQqrYsIAqCVhWrnN7erxLeY9N3w1
1wydyzCKYFXoQAI0JtkfeFAh68Hnya/zJM8tYPiN7FOX7m96ZS1ofWjpvX98vPYM
WQFKb91LIwOLyvssSeQVPMswMN+hl+R3GhZFHQqh8f92nkDJBXzFsldcSk0O6Vcz
NGLgLIMWnFGumldjVl3t5MqvCIZJ7RyFmHtRRUcewZOvpyHuHuquvK240TQEh6dh
8Qp+tsmTnrRcCIAIkFtTg8wToM6/+y2Y5k8L9ZC2owL0jo7QusHgxrz4dmaf3Jim
yLYPXcOLEnCfXLu5hRhs1tJTfwTxJqkPgdtrI531XPLkFyX7Su2L6SC/73yaxZ2y
zlk1iM3ZVRL0pl/UKsaFxk87jhFyRpFKRQznSaXsHrcIWEGh6vZWWBJx5+3Fho2c
plKi9Sc1a1qBc2uRfVEoYJU51cvy5g2rcD2R/Ilsp6WE0N8NmmridJSN1jt5qG0a
R/0OfXVT4qkfb3KGrQF4v4Pe3CJGsaiClCcqXZZzkxc8onsclBgSroJF/h9LDAwF
YxBS7Gl/HSUts64Ek0+zUERM6GdyIuUy/AGvvKjmvT5kbKpi4klMddozDtG/MV/8
7cCRhqL7WoZId8RrWtsrxacvSPdejWLvTRdPAF4FxIxypD4Sun12ZSd61x4XVGtJ
iC1ceSzwzNNunBhHZ8gkPzLsnC77z+sargqINxueGZ4IDOZqpB/G2GyCJGroC7JV
/gZnyTXXqpb4D4lB0cPyPUtfQbLxO+M7/4LZXNu4CHph6yxOlnaX3TrV5YA5aBO7
wpxId5kCVphNHWzQMUzrjq5WDRLYQjRwkP+444LLZSgLc9UOJb+lirCPhZNKLrlU
fnFjLieXa7JdVIU5oXdXzpkl2Sx5Tx4BFoeUm0AnJqqWkuTvsVOGpo+yv4PTLxMB
QpCbMx6Gwy7M+94/NyCij4vyQy5G1MZPowNaffoj6DwJvBheKvBvynYbsXrXH6N9
T0eIn9KNAG1Eg2xGtFxfCdXpXlR4ogjMaG6yJZ2oMqQRoFfhZ6J0i6//n8g/rpZj
mSohh6+9ztyV4KD6b+QKi9swVvPCXn9WASJicUjTNFE1QCII5AgLYRasL2ew++TS
Z+mLxbK6xETmJA9wXvyYl5TZpfnctEO6OYsyp5ruP2U8+I/ZjsF6nXJgU7UZMv/q
nW1Ag6G++2yiH2gTCWzo28wrGeYk8RKeGXX4a50kvKaBeP25jt5eLjN/5MC76GJT
g30i05ol9DFCKxWEnSbmAk1rqsYtZEM8af9rRqjsbeBYojrV5gWEoZz7xrTnFzso
2AfYoq1ak42wujJH28RjgVFh4hDPIXDqpY5iuDqEz50I2x95S1SgaUYRwLNYP2r8
mJvIVsmNwyIqleIfQKRTkdHJ9oIl9nghTvu9J+bHYURvxqbSKSNsUfKEjIH0K+PQ
2nqX+LCUuiVun8NcUrShAxe1sXvZd0rDU/GHgHm9SfDys1bLxgo7s/glaGKLy3bc
ZnykfQhqk+XK0iQYj+P7hapt1kM0/zavwVtHSlwWpb3niq0wMj7Tu07+t3Yn0raX
kShurzMVJKBoevIma4PcjCRwiEoxK2Q7gOMrA/PJuCyd4EDaOJLZPb2lmjdDfXGJ
r4cL7CXJ01zvhgWKTVGkpYAE5/iJ9KptNLz26BTVQK2XoR74zfOUhbtWh2jQT+Zr
RjVoREs6eq23zqStK2A+qDTbKeZDvt92AyVFlZcvYjt2su8Lq7itjmZWI2lmosNv
bMwO6Zu6tFs932p+g6AK+ZrM69f0kt/ij4SDBM8AL6G1z7sjwmTPsjB400UF6FBl
ejQFEr7O3m4SH+j2Fxwh74lELg/pN+CGRfyBffFsGtq767/jafuESldVYu2l+wSD
roaystTtNQFlNBEDwizulZDX6LfZ6ZcKC2Nr7lAXVFcCzj3hL86qMxbearERW2Km
4VjcANLaiZKYtoSWwG3EZf9o7wE55+enSdjX17ijz/9Roc41lwGnH2bepELHoO7l
Z6/y93CQraZj3iMmsjYGxLBSwlZlHrt05Z77VY85K13nGW9Q8xW0bQm4tnkuDNid
DqnEOKGV0iiQiXm9EhfC/wdFi/63o5rpNXwEvePZLt/tTxfyFAFlYJasYb7zxsU0
vhFrE4tgnY6vryYAfxI8wuAvoRcw1PLVXRO25h0DymHLhc2N002fV0d+cP74ehmu
xle6RbyyoiMwOov9jppv4j9An25/Ki5cOQAw9HGGoC4Jcn2ftNmwPrbK+8WMaPvG
1vUTzsF4u3tcZVqQT3yVPrpdpJmoW3fcWuqc3mN6X/fxfEeP0xJ988Wr/Jrvj4I0
CuWIrYkHIcE8SGUPGeQwxmsS6lVcpJA+bBoxAilMeQRHWwSLRbRvWH1UrjDiy2zS
JeP9TFBNp1+unV2CaNhTQ62TnZGd5J13CLFYWD2nr3ASa0v5OzpjMNf1sfiR/bUi
YJ1lgnrqjy+Mc7Mrc2Bh5TEHyglUPFkcbhmI4CVwiquu5JPJrPrDrr7sljWW1gvC
ybXBCNVBh2Bg5b/1h3QxTEpPFAfZjAJ6+VOL35wpTN2ZzJ1Qi8BXg7ViQkHuty+a
e+9fVapTphY6j5B2IoB0kLEVMN9NSHcYUFNw4hssQ3BbtZ0faL28GarGS/vRoKGi
AHuALF7kGglsEBpZlbs5C58tBJil+pbfHps/HWLc1vGI4TZFR88GjVA3asuj/ya0
LS6IZQoV0bMtaNyuaEiS/tnqIYlztvNxbQlyTIza0c4EzAXl0XLK97W3zKvMnuUF
ADGlDEs3LBec02F9m0d2+5qu0dQYboX7WzK9i/TQq+wQK461lyRFtFrImpI6CLFW
lk06HHEznAmLIMiLu/IdVAbHzr7PhrmZCGk7//+79uVtE5EKzJOEeh4Wkg7K1z+n
Bg+tPhAV74uzyEPsS20QcveEwUmq0ZVmxpCg4UngAU6kueimg7Ex1mpEDBHPdAuD
sEQ0dw4550hutj6N1lKYkpU2JfeN4Qy4aFoy32erFlGaqXmVaKl0dWjoDZC+sNST
5uO/IzaeKFJw22g0h/X6AmzhRkMe3jDLbVmWIqbUlswZj16NGTSfXAsQu0JrmLuC
ohU+t5MTpgciBNPxh/WwCgbX1fGYs7ehqfKdu4iK6UsigG2EdZSKREosyBzTON/Z
SDv0Jc9fo9UVVXMrNbQK8Qz2gh7tKjTILPf/D4WZXpcofz7aJgLJI4kCJlhch72p
GOq1MfvGifY+haea5+aR4IWTZ6hQ8aS3PRuEtmrZz8u1x2EKiyX4oNPM/X+r2tE5
cF0A+ppyj5wPuQGiZlfBHz9AslXKiEMkjTP54sVrzGB0bPVWNS3cFK91csBamlMc
L40XU1OVfY8jbKYXTr36R/Tk8JI3oQ9MmohDPgmDtqUh7iGo1PwdyFb/43Y2WhV1
2yljO81ZbW/zBnBHPY26sc8yBb2Re2CoT7amFoIqzcdkOgybeal3UKF8ghxZ029A
zW7ZMR+y8LoKwA1MkOmYSlgdXz4zVZgbevI3VXeAH2nFez8nenC4t4YDSS8MWJLy
YAqw4Q6TczMeucaq9JojQA+MURU72Ls5bv/BG9Ex0w9dH0aod/orzRELVsGePBb/
gdNq8Ay/1DGUtGMzm8QgLdOfqffo5JY2TRVr3CVnJ3fpY7DHqdxq4XFYJB1ZpQlC
YfxaqznKIFL2MbwUljNlFGrc1fgBlP7ZLMQr96UdqYYppTJB1gq1idvy85Y87RuV
UsVHuw+IP7pETiyY81Nfiyro7erd5ROx+YSwnbxfBMSnIIK1VfpiWVpOZ3cyRrAU
LsqbqCVi0tbtjgqU/7b5UUR9Y0YPwBWs0tlodd9dB7jxx6sXj3apYkul+We3HjW9
6nM4u9+NEvk2SD86AhpE6kI0r+K2Y3qVxAD7GDTUxYI5md1t6cRmQDKU09+eztCi
z3h9m7ATQX0zmc6E1xvJUZfYocmBnMh0HKCuNGkDVBNCyWCPpKWGEFxwaMCdIQSV
nI6uET2Ll3dCO5GKqZO+BqI0hXjy5o1VQf7IvBMGvtq5zsEUWl24PlL/lyHqm69f
+OfabyGu7PcrZM6HQdUB/wcVy4TLP0A1JGMQt95OCeYA/qR+25B2Se+m9cJSD7a2
GD8oWkos/l0hAe3//wHHw1SYwfJYBj/8DAdl5pwzUUYdT5QDgoGyiI0UKNcTgDD1
dohp0m1s0FArOwRC7MrXWrI0lL9dXD0ee94bY1cweUyYExpOmWNuf0+7u9s9+XCa
2lXatQ2JT8pIwDo1PBnVNwtUUvzMfbGg11LW12O+hlZmcv7Uwdji/sUUF/4Hp35d
W36FhmpG2Ayt/PjClBOJhna2ZqvEkTd/T9sa/fO3isXe9Un2CWwBQZkvffqhvkGg
uaV9UKRSSSDg2CYteuMFh4nuOxVVC77M1Pz0u8I8Kd6OrnNfn2e/6R4280nrR/kW
krnC3H6jUBQSRUSvKkmrZZS4/M6qzAcPvydbMhdtqb/+uySN1RGLxTOfgPCvq7qB
GTSJoHEF5Nl8YvG5KM0I56ILL6KPn+Q1AOBz+QS+IVoehXyfuG88GMH/7bIKCnoP
y1NejNycRa9sOdgCfWWUL8v4sypjJYFikxjbr63B8bf+zIOkDN4ifrcn5Co/I3N2
9CF7/8YWHqS8zIek3vVfHXOXGlu/7MYiaXDnRZMWR2x+2W3ZDOkLNEy8ScyqZpMU
atb5w84H3prFpf31cfZEFkLR/89ZX70NJuy7/0ufCwQW/e87dPCHQ/n3nL9QBPto
gHdkCOrSaEf6i+Q6L1TIB9FvRoSbnnM89v8/nb2N1MPFTcBgZ/cE/rHxsCSw5wIX
Mr1zXkJ4KN/AyohjOSahBsDAPYo2lbI3BVmwYb4jvKPoiTpoqtwrwGQbVnE3WIbh
xjkO7+gzHH0luls6vkD2SJrmaPWyqhp2s6q6jqxl4gp+sBux3ccWCu1SyxKvSCSN
1jGl4Tpgfpjy3cLkuAz2/dlhQ69CIiSHA4ZYf62k0Be45UcJCnCayPck44PMiyD/
TvOJ0AH7x5cG/jrd5PwGZRBjNsnSLMYcOhvVPxonmBqua+hqKxb5p1sWK9WpZVyT
0/OBHqu61BHwJlyMyixrW1yBIUqkX98iOwsWcEjkjo+TnfDpd4TBiUFt2VsGUxau
CTYCSmWva2I1E0m5B+SvuR8LPlA5Atm5lLGrDLpmOKU4L84VLfoc/RRX1V6YEOm5
kdf8c1QlFbEhWwljds98ijdhy9U/122FjJeyY5kx9TKBFzcNyR9dd3BSDy0eNj1W
C8py/z4h53H9pHFbUKR8g8zySWSb2lTfREP8dNb+Nss8joIuXLr2tEiWk4w82MIe
KqgNp0zA8wRKKUnuCr9+jpd2VFZ3Hd1HeH1WTNr2casRYYav62OH9iwklfb/B9eH
V9pCd1okvl01Jy2Mk9k1MM6IELf1HL2+dxJtn+q4AeyjGXjyms9u9app6DW9Kj3C
SZvlZlFwiF/sthfe6fBB90qJRzpY6vjUOb+f9lM9X5DLV4hrmxeZ9D8WLAaFmkC9
KAdDmV5LMDHNJbrpOV46I4Tr507mG8YZZ9p8kwiizZ7U/uJOJNZ5JA4ga+BcQmQg
nCqATnYRm0yIAbzgMv7oDtWAOA+CP/Z+eh8huz+YIZ5wtaePaabusaQ2r/zVdwWL
rM6lLW4m/CZx/aaen6Ftky33c2oge6f3Zre4b9yn7MUA5XHSSrOI8RJj7w8ozmnr
Tp08jbcI3o9iXt6qqCNJLE2tOHlhv7cpN4zW/xAaewAeV/urU7se7P+wQMIANRdF
YkdPvmuxK+3Hh2d/AhbI2c+iYJG4WwlfzV9R0esnE+CUkWtVPVA7V/W9VHlo9CfO
Vhf7/kLP7kQX6x/TukcO2D19zIFv2NbZJeDmqdb/UZb/4xtzKVR3SayDjXSpXAYy
ywDiQJZURDc6H+r8uUXs3Viu7l8s6jXMtlaEwJPW4NakpD11A76aNlHfL5L4PXZs
8q44hMmWEcX6i+ISH3SjLogDuTK4OHDqg+At/izVVu2FxgguOahgrmsjPPndA7rK
lCws7xf1U5nV5qkfx9IekguTfZvnC/xOgcAW208Yh/q8uyzmbbaJscHbrcDPQnGm
hAfUdr4Dl8/vBn3FU0qO21DO+9bqX7LF9NmvIWnZxP2MyMiUG8IsFLhwuAY9pZxu
9I3OZ9w5XT9mPy6Fkbn88lEK8RoS525WFq7kFeM/rX4xrQpuCC18G9s83djBvR9w
NuGIRxOetoQgeNgYIvyvtc8kMRlrBeL7TUcjeEQKw4rrNteKm8DlKeNlPN7A5IFi
7mvgFsVtQQ6N9HtRbuwKL1xBd1niE1QQZXLYC+JUiFGNnRlVZPa+PKrdX7wK/1MG
0Db4viwDhU6gVj+OAkQnx5HgE8fcVf4k6pgAIdt4M8zciNaZ6gMy1DhKGMc3cB0Q
uHXFuKxsRAcA8/urvAg+48FS8mIscvRtYrZPZ8JI7KMunyUiCXchCjiNqLGfrme+
P4MKY8VYVu9RfhS5u37HH/5zZ4KHkoFqCfYP3BWxh+lCKw6+6egrnJzoxofzC4Dq
opRlwnL3+JUWjkMkGBVu/5TgmlBuc0YWjn2Ug34PaMSGWXbrI3KxAksvqRDQJ9QT
E6bI6XeWeGb/MQYKTshxlKrpBA6/nBjuKZ1zoKqwzBZgy8AaZJ2JpUaMBwqioEgP
8kYqGx5iOg3etXBwUzHYtadhB4wCIc3ublfenQwdEKZyy1pnVFtwLaZU4anhfyyD
iKrpk3dM3+TkTimEEhnN6L8NaQ64qx+YaBIdNFuQzFNJ/3RvvB3oz5VCL7fy3u4Y
xGjXqfppL0eJ5310kKLuxnG+MiOpdTxnzbH5B5P4szIRRldnGQOEbIm7DQo4qwQq
zqJeUrFACunlyN19670boPBclRRXHX6kNyhoxJZKdaAr4yRNNsG9VoXZtOL5YBVX
Nyrtj1GTbsmOKMF6oevpQGMY6dBhgq4WHxWhZFdLEJQMsYfNzhglbmkHJ6nszTyu
3MvenLQ8GTPFIoWmt4U/W72fe+YbK85tx35qhjVD72lRNczknPoTUdxHftNGFGts
OVmmHcFe7kG4CyoESK3RUhDu5OUlgj8F89gDzGmDcMPSUjCw16CqDuzxg1PeJ92L
EeSNUDqMsI/aWx3nGjqceWcc8lqeqLQiFhQoa/OEvyYG+CfI+1MmTmxeagYv6qUA
lcqkL0LEtGsD+PQGtr3UOdKlKjqJPpsgv3RXVgy7StJGekbbNCSRjI6M6fRM1zCx
V9ejp6cHQRMGwe6LE3cXLEm8Ftr26Y1KgN9nm+t3lNNR9QXs3YeZtCKZvWKf4t6q
XSNCL+Q53q3Aas43kY8VD2qCLGxJYVXe/MeDGPhBfQa1poDzKPrn1jigxc2z+/o5
qV/QYvQee5V7t5ZESjqQkrkca6yyaHpAeRsLgJdgBhjjeG5eIN5JJoEIvy2TOKfn
ZmAk/K8I6mYb+UWaxeiRmFxKF8HkUZTe2+rrqKN2a8DqDry3t5UFemINMZkWB54J
mg7snaAknZHHw77n7jGnd+N9sspV8fiF/aXVNQpT7qesjuZp3RZ13tFAKV+LP/Ev
2Ch9GuRor//b7RLNQO6dKD27jKncNDRd5Cxk6RctCReDGcAKdDArGz+p80zaRT1i
dNLgIT5xjtRZwQdAKCKy2UsH15ktcovjgAMjTdk8cRfuX9FTgjgxhf2yoVB8BgYd
o0PX7U7WxTP1j8eOugABwksdaeIGLUYBFdcFTSUdE1wDCaixNNqeoiJP/93qxQPd
blnENKhm+IzOyXcHs4CWHU0MbEEg2/ZhpgdS/H6L99bNBGJtlPps/hVqzQ1HA11d
03vtiNxmem7GhT6ccCeOJaHiHAhfNij6SUsmqN1nnfPNw/CSNSVYVK3xgsegdYo0
koyJSoiTu0O59YwLI4ik2mVziscbxTvcxlfrXgLqgUla9uLT0KxS3sd1VlIqRez3
UbwGK0vIPUV4COgBBVnNeER1fJxkw1LP0DJFJI10s9FXTYZIyfhtxFS4PGx64lL4
ssL1VzEcqLxg35gz2lE9TSI9iNNRVhlfIqs1MkTIM3qz58I+iGbaM4mJASdd+uxQ
bdhEO/YcaIfyXpqIkmdCGidLZBqPnKS3CBzzr8XZLFnOHEmxdOuvIonywDhSQUh7
Vn0lgMnAEVPI0xzkK7S2zm4trM2d+Ggc/b9shhGSzV+rDzaj84kxJst8ZOC3LOZG
FlO8nEZIS08KHfh8U9ysE2aLlqofIIbJSvycuWBugb9GZNi8VDH4aoYy9ZijyugL
q/SbNRjNyuFvl3bLMNO7+X11zqNjB6cDJp/2T1uTznnG2CeHAKneSfhLy0d44nlG
IuODgJhpOKXDZqii5eBcn03cDflIhwguHP0A72RI4EGf5TLLadffjNcpOFUPjfK+
XP+rFCTi7V9S8NBnyxI4tZrK+tD4MclQ4w9TLTJ7TxHkxfkhsl5GDRsT0auU3+IH
FR7fI4UlaOSYxIZTfpo1bsS012JvZpjy99W9T53WkbqumWn+VGmJGB/dylhw/ZBW
thfelMTCfTtB2keMmORBM0IUcSprJLJuJH0R2brwKw62I0CFUyjVti+GC/XWZiGD
dWRd8nOp0GTFCtq+9PHGrbyt3rTSFMV4Kmq8GJlHAu4c6vb8IYt0cBquYAqSrjrl
syp5Afz21Q1V+93M7IPr/C44ZpKgw5QDYa6FieghYUQElbLGFuU29TzFoWqDjy9w
x6bvKvchu4Yf388AyScJ5BBtymsGwBHkABffGGEC08L8C6tujFkzeGbWfPM72WWt
H5uCVEK1W5NW/BkchCK3sfuyiS2AOu1TKXjaPkTngABszSl9CqfTKw0IqxkdgNBA
0coNFM6OIfNQktSlT4rcjwnSP2scToP8RwN8E5Bgnk/+zNEO4/yEJzzPu/lgiFsL
r5tfA43WiBlTVTL92QC5OR0qsKHIBX2Rqz5Gi/CuwK1LKcYgf3jFmLW7LjX6xmv6
CqOInAvQxYsJKvreQXdxOVRYRHswPWHMk+4k5SANTYib3InPlmYrkxPtKmqBiaUf
SXw7Of9R4Vf9oywI9Im5xGZwFWTqnSOn+xv1IQGASe2KLaOa5QIOHRiaKSK+7eeu
rXj2Vbmb+CFClIVLEnsAtYS4mOESxF+xz/KCh4zxTUc3CBROztZc7vlY4r0TSVeh
IUhkRCUABXsY+ENZ5CGAIXeADpeji1peK7JqhklP485cyLPg8qtW+9BnTlVuNdzy
YYHi9Mecvrz7rCLEtDjtcJANpIrJN7DRORXllYiHFmlKhBJLycTbVYWCzt+ga5J5
xjZimbltcOdVFcKxxtYjR6cyiapnYlPnfWpAmz1llq+c39Qgl4O5ENBcbt8tu6WC
+Mf9BoTju+6t+b54MykdIeBAc0c66Hxt3/gF+Mk+eHPbhsCJEipoJLZ0NZd/+cQR
sXojtqOKLwUq0j6SmMeksIiB/bNBU6IqltQFgC/PljMpi/fCeDTO3rimyUfnx+IT
vzpLSgAvbjBmGnlgXVmIdFg2S+2weV4vMT0Bguwd8re44cjm8t71yGHQyMqvP2SO
OuqEtaK66Cp+y8Wsj9dZ3GSBXlN+ByOLlYGCY/MEbvdAE7Ci84tTzVhyRE3X1fZf
nSBwDlnoPU2nuCeHtIB9aZIa88TZrDenPPRHwCQxQjtYIVMLO14BX+wAi2+j60cD
qirPFg7rQM2kv/dNjbZs3eKJSFNw1Sj4+sYWOmLyOhtJvz7Mr7sBtTsu5THqBHM2
rlsJ24NyvGgZHxUpd1V4EYhHWYlqB1Bn/pAn6xPB9yvZLlj6Voivt61hNKWyiO0N
wNFR2VOY07vlGnRb0MxXCFCdsRufi85z8KlBBwrnZJHJg6/79V0zCisnM8tFe7CT
Iqk8CCn7XC0MQalUOIrSLOCr+5w3z6EsOtbG8yXDChpgIOg5Bpk5JXOI2ugsjEaC
73WWe6vuglmvcksYv9C1ecg6y0Av4YAPLcUfTiktPOy2ERyNMT111PbPiCV9P/Ah
ctypQ/DWTNvArp9PvV3RrIWlAueEsqw4ocW24l9shYkiqLhDmUPRmIVmAhgH7Rkq
ob56GReMRqFtkbfKe70XlsIY6TpeHSyriAyGl4iYptdVskfCoxROnPP7GHBdJaSw
/cBAKckc0Gz/r05Ds6N8UFFZecj9cIKQhw/1ebwtSk476bcfALNI4dtBfiDx/Mkv
HsaJCxH9evT6FBBjyet9SbgKof38DU5JAq2vQFuEqxlkaoASf75jJbd4hz6JC+aF
0XxRIS7vDCeaZHXCIos7F2gjJnD5vDvWf7lM7Ayu6gNUL+zxDPD/DYWdQ4qHt8jy
dIGdP7OVAaw3YdaVGhIvvnmQuVms7gPqpw1o2/Q6N7QMNB63/XNxChVW36mInr6E
INACQDlLwoCJkuYefr6Xh4svbTd4WTwH5vCnfDNwcCkkx0V/DlIMA2tdK2NM96B1
MSSOdmDl+PgF5qL77zid4Twy/If0lhco9mEHYR2mwWmpmnHcGnpksu+NCkeSjmDI
mdCCnznimjo7yo7kDkIHXvhMyx6MwlQiMOFO0ecxCVYcDG541642auSPZTo+fjvT
YaOehiWC4r1ZHaIJ85fcyXzYT3aS+J4zItwq9rsg4E4UfN+JvekbqPWSxx9vrcpN
q+UX+zKlNWbx1TKnqafFgPwaCSc42gju28+yPd6sEA2HgUVd8prFZH5sJh8zO8ls
t0gkosvf0Q9xi9NwwRpbyoR+VK86FB3qdyXUmDwJfsCq84omKGbpACvNl881npfo
oDzbYgrQyWPnlMT3eWImO6onMfH/dX8L1g40P0kdN5M0DhXMF+8N/UP76tGP9uFL
mbSVxlnG/Syu8l1XoZXq5suPnfMlblYfe2WK1M0YzywgFetJPRfF1Jved6AIquFO
UMtuX/+uFGe4x+jih3SE3cuOEszueZsNrn2l5qDn/dieRuD6cH38/BRJhdFsn1ri
TnehSOeivUyZflhnn9cxxRqBn+55x96oNTysdglW4+HBCEKO9U/LASo3czrpE/RY
BTHNlCxevjq0bSRk+S4qA/f8zz0p1EF/WbeyMuVqNinv3foo+TCH+mXv1UCuDeuC
a8iwHld/ZiekkIiFAsbmh6OfVu0khEMMBZd+40ZMwpAWklsUNSQNb12prnnUf6Db
9wWGFhXSzNLqPMZXjBCHdWzn+7NNIQf7GapAjKSfxb+l9utkkQnWx3jMcAefYVBs
l3UA9XRbABQwaGyreqxn9DSklQ4WzEnoP/d6jEv0woBqoG7dAhFm1AZfUUpiyqsw
88+2pC6n6YHqDdqwSIujbiyeIn8YEE0VJhDP2FHGjs7wF7UT6+glH1yjzduoFQQb
NwD0XdsRNvp8W3KdbrkYVq/zlyUhEEMaF70zGoKeujFGFKWfZzCtagoyNuNmawSU
5lsHR3XLPiX9O82i5gecUnMR+SBUVRJGQFzR8GRikeL6w5UedlxjeQJtQOx9TAiq
nmLmNhhD5Cg+a4sGlUL0IJa284LlcrWkhbu1aLPF/nYrNaEHSfhiyY8PRFXQZ6WB
06MAF3OiiWGNs1pmEAyNHzc5C7ku2PBU5vKYb4+JKUwva7RrS2IHfutBJttVvw/Q
dOTvRS2YWPrCEtgUNZEPw3R96tEac5uv0ypMJJreEirg3SCiGTGgu2pHmpKDTs1U
eJLZXMKdvV9MdJHcHte+woUtWuKscCmDX6hoprMoBM6C0EPMBraVJl9MY6f1pL8u
qXYr4SRqVW001WZBSM5txREFLLM9223tARJIFN6EEsAhFW80Ds1b9cBEhnHhK1QA
lGTRYT521/nfQCiNc7fMuiBbVFEAORgiSAeL8W3idij89WIMSRmjzCDxl+ZzxzpH
IhQ+hwWvcKix1rW1aZ+iIGmkfVib4qHigOZ51bhIvkby3+qXx5oi6q/udEZG5VkY
2JHO/jqaoTjJaYaGd11o3HL+IFY5FeYJHrKOW0anGNFv1WGnyjXIjOUuQ4pTT4W7
69yG/S/ZynM3GZaKl5Yn9A+3PhNwHg3oiHbjNMIV9CzB8/EWn38biavmQgfmNY3S
KPA8Ox4hgr5vx1VgCn91uXvaUHS65LEz3tlEAOiP+53QTlGypbky0f8Mj/G23VxC
dZv/ISjA+Mw8gg+6+z2GOb2Q2tIcHD/SGi7K21Hz7RsRjgmqMLSKeysgX0WLQPZ0
/uBgDHwYcMniCF0h+8O5gnb6p+b4+Wn5TQVHmZ05BS3mgfhdIhW/kgbmuTojaDK1
t2wCztd4t3Or1L+uHzagpaCj4sEZ4LYkXvmfTj3/puQu+y/6OaMUZvpzw2psXTHa
8WqZc+ZGZPZcf59TeOZyvzFgdMBk+RrTzqSrKhPpUlJfcq+Pub26jE/+V2lFMMq8
M8ekeaYtHPK9hwmLvN2efkb/LoSZOQLAYU6dsslTH1DcVXJm32BMa3I7RePHFcIo
exU6ZbPEkzLheHxflCv9n+d5Weq7XIzVBLU7Rf05T7m61SSdmxs6dFRvnQph+yjW
I05jJ521a8GHFO6oiDcJkrvbkpZ4QBLPuEloJn4ioYRsS5em0OFkQGmyrHKCX6qI
zhl+dvIC0kf81C6eVJcznemw2Fdy2kUU6gQaE5lU9QN0VwXwjsGnjHx3nMgvlF+C
FDJ34gattM3eyFpvnKopt7HakQJf69A72mGlNM0HKIdvAY+K7Ck7VAJMa47xRshZ
zHfsw8T18vcG6ydGbAjfUIjY2rZF6I7qHi3/T7Z/1VgMssqeX2CReL/BVyPGOHBZ
g9ESTAKfCke2/ju9SAVJJyDkfGOaw3pRY398lgSAOp5DoMke/w1eaUMBrCaCbt2T
ajiOKJRiRowGuOX9gWC6/Zi9gTbmuPfTCNhDujfpPnbkuNcp9w+3zLdSPpQQ3J59
/Yv0T/cqiUGTiyCqfvsKob4tSBH20xajkGQMDkefEv1szC9mDgdsKY8+5P2vMP/x
lGuSDJ5IRO3F8EJN3JZgNQwsC+tt64Ja/SS+/zVMqc7eoWFxyoGmvzlWhDsD27Zk
g5un0zCdBEPp6jfgsL4utC8H1eFvQJbYPfa/4omcKxudK3QltbEwxhHKpnlj2xrC
ipMgXcbaT9+zKYVlDbWhk9CDvUZ9pdA/u9ZRZNlZbiwMZdivML2aG60sk4rwRvCk
mu9Zbj/289iVADYyyrf3wmXutTarhdY0APdMB7Pi7X0gkrqc51ZR0IlYSMJw765B
J9yR1l7KlMinUuZP4QEGRYWnZVhLho0kXYZdLj29kebKQxCh/utpeWfABisFFlgX
OsmLxRMkl51DuhBRSVz4i7OMzbr0ZwSVihRmL459l+ei82LnptfpdeBZ2Qv20yhd
Te1XeHBumkCLcBs0rO0naqvzD63P+z5G6OttJtkDKfJCwUzBoD3M5uKk9QNzHTLp
EHcMVpojYHoM2VgYXHHUj9aDQxa2dpaNgsKWGmzu5YGUMghCo0Ri49OXnFWI8RNP
vb54J4t+o8mb7SqPZgFiB5lzUFE5FrP5SKKlXsXvF4/tMX0ebk8gFPE+lpxNdnk8
NE2iAgr4ouE1OWqiKlsdO4nx6wPuUAcG9S4u+gaGueCR7ydgUMngMJ0B1BDbPZzH
B7EK+hMqWGgAe9ydvOJ05wfwvU7b0WjMC4uv2hYOd1qggOuTwY5S+vRHMOmWuuKA
KD8rjyxKBf8Lj88aO+BAjvqLlFad0ky1AC+ihZTn0qe4Wbxo++Ow5DDKUnMCWJ0/
lASVOlhTRz9a8/nvVuhjZDYcarqkJ9WottjNKbjdqbncu/vB+KIpE5HrvdSwdqhl
Xrlu66QdxHST7KLhXvhhatniEmV3GYDnHG05mEgFvQDltqeLbmdET7JfAXqjc9Y2
c7IyLavhXzEK6HdvKUIQ5exi7k9EEEqfVuDT4dsIFZY9ubL4+5qUfjmK7UzDEFtB
eL/fIOVFFmji7bLgizLok1QIDjNPrzt5vUdUEqe9TCIap7FHygDLdWafEJMTJHdg
W9HrLeo7wFK49iiXFeHKjWePvu37JxWE85sLSIGbfEpUnWeT2tZ+MHtUqnAKyhlx
q+hC9ErUWeqqh8U5cTsHn0J7brK6s279Bqpknht26MxYp0JuIn/iQqFuojEg68+O
pt/D4MSI8BLjEO5YbRp8k4yv5MoR0rgXwK7tevMDRBV4O/+PP78mEbR2JXuPfByZ
fLFsYSAv3K3bFIFenKwPRpWle/4ByWMH4LLBybudV886HgevefYDiTycOkGAvz/r
9be1gAmZaut2RmVpvHTdh9ocKi/y6Qx/UuqoUQQnuyRqeiBNS6CnGLJt6TXL+BdU
aj+Wnf6pp7dHWIinEwJK3P1heNvRsZVE/0kEwilSACcg6ZC37UrrqCYjOrf5J8GJ
o6PrwVkvzrDCpVV+bVo33ck6C0jLhfBZA1Kh7PAoZqXMbPx5xFIux1flCeRPrl2U
hteTr97BiQO4uGN28JsjhCnNSOeSAC6aMlqPsV66BMAtG9SX+f/ilzOEtTB9UhI4
NULn8J/mjx07mE1MoRf9/F4l6QiuzPFl8huQ4Znk06a9+qXhTOVm5aGVd+o7OgWe
DpbPf976YW6/AGM2QLhTwFNBpbc00pfrXKrYzJkLjlxeR/iJoftHmFW7VakfmIKE
/JTJZIWdiPVTIcCAjCPlfgXQfldwuku0o3EqMjpkCLN/a/vXxD+Aeno/luiexDXH
zbP5octe0r994XZMYeG7xNwfpINYgMKed26DZjNJcKi9fdlbYWETa8bKwsvhuueA
RJ7E6E7dUIwvraEji1nQ5kOHpOrcvuekW7e1imlGhcncdysnDi8k/0nI7cHfcomn
ZWLdFILCNFUqhkJwso41xl1WQglGl0sCXBvp6zzJobuWE/7mT6HcIiIKfYOAhT/l
n4vZj4+9QKTtP+B0XYWd9eut/FfELisyBGE2vORMdDM4aOXRyP683Kg2f4XTeZfe
RWzCURXt0GMuvnXiK/V959An0yQSbJ479F8KYzv7ynAFel28Otur1NndOgYnGrhc
6qMvVUvPVLRjRehM9N8WfmX2090xbJDUy7D4yJF9dmWqyHxT/KDnRr2pFlz1yj0f
Z7DFhA4G17CWwgl0YSLjxtrDwaoxgcUvLWDOYoDP17y5Fn0nXZPWNtCjWpDoRR4j
2VCYjhFGabg9K+qPWHYnWuAW1mMe6m/7X2dGr5FZrvJh0k/AUFa+rJ0BY4DnqikK
489T4Ga0b1z3pdIuvt4HYvdfcpzBgFLvZMIMwOTMgBViAhofnvqiXsO7anSK1r26
sEpj0XzW0MTki7E7O3Kozauqr94ZFt/YqKyERAbl3dhA3TZ/3EjwAX5tl8phNfHp
+UL3zcPmLnWu+/3wRN1kyEpttVpDXcOrvwgxb10ysArhS8+BxJ9iR/1BLkg++T2j
F3OcFkUtE/gnredZRI71rmVq2rTChPDWSuN3kn7j1/cXqgq/d96ytZRGe1YIKfhz
w+GsNu3GOHYPFaebDvAqwR4+Q++MlIZW/BGf1Qn5n6/lXRa6dn29EcpQauVwftKX
YXjcwxzw5NqpNA4htRSJu6Q4jeLrPSoXNNWGRZwqLYXtA7HTz+RxA1ikXCJxuTdk
1m4jRav9DOv60wVipbSNhEQ6PspL4sST+gDCop5DJ/7G6Ai3pUZq/Xj82MnGrPTB
UNHpaLH1YWME/WrJ1EX/Kg/dNpdPQw7CRcm4yCVJIWfw2kTlq6uSRs/u2A7bruIk
Rvd5UxQmPpyp8vX3plJruunoH6AVPlIhsJxttQlXrcyEkGWChgqN8pEeys+vJoQ+
HGOIVu6jA9hoCsmaNeCIe2jWw3oKRRZ7WNXFTgNN46UGHlKfJXX2sEIF/6m2kfKO
Q+PnWt5fOiJ0SSlXCg1sS4eSzEFPoFghHZO5atzUSOcjPzCQsFeLot1yu8wu3Ynb
vhezAOmT+eccsLK/PDAgUkn4i+ehtnoRv7f0ZW5pOng9xGY3EIBKpcDVvVS0LtEU
BFYyJWtlHgVgQ8qCu0TFILJqiKvVd/sFXBsS0AQjuKIP3NWYpBQMrAceU2o9ddm0
K79qkuoH5X6rnH164QwzqAW7beQoc9TjtBm0HdaHi2nSTShr0qlNI1FiACLe/UhR
RulFNx/TtfzHOiKatvc1u4CsQBn3f/3so1Ul3ztXeGnnVHoX833ZtlopPHjxMl30
Xk5h35c52ZytweJ4OSW1HqEhalwCYsKeNuR5f4kHJxk+ZuJmho6/eX0N7w8pzA8X
P7ba1lSJrn5oPg2ra4JagN7bSjDb647sXLCfQSrN6/Znm+NBXyxe+WMnCEmMHBtM
K6O3XDih4fY2KXkhTcjLJt1JE/tr8PIUUqBtPhUd9rsBy2XHIgom2Dt7Reyhr6DE
mwq0jvbYyOcs8b1XG35mEhTh7eb7Mls4feO8uEaulreHEiDMxBzdwMsCJWC0k8YP
IcFXN6FDyDP0YBWsSVZUiTH7y8qyZglY1Eo/q+xv7G8ndwr/Nnlhl5A6JZ2rqoLl
cdmvgmQDOhH3DmIrKY4S4OIfhszkrky1FbDxYR6Pe/pTx4CQwbVzw2wTD64xKULa
I6+2DaV7xkKO+XmM++5CUKbYI3e46bRft+ash6Vn4JiwsWWpYsd0XD2pZs+0hxLG
xFWn8B5ds0UCUPFooKu9P7tkaNGCGNGn3/XKy4EkCqJMV2ArFCSM2YL8rX9mjlXO
wIvAfC7q5B8inY1ED/QWqtfpRR944M8uRGhlaCzRvIYqY8NIYg7pOnD/1IoTNpCr
Cq9wEdEW402Zd0uHKJQxkyTLwiCqrQH+aKbyahbsb1U2xsO7ZYMhR13YsnMAS251
tIfXVc9zM5vLBW71SMKjP6P4nDxtTcqYdUisqzUno6Ae+Fp8n0WtnEg6o71aPWvz
T3sWDx6FhEew/T+cehDHQJlgSAQRKAGmyB2i2m73NmWPWVLkoi+Qw93BAmzLhhtc
Xrlkj3uCeAV2HkksNMV2HvpPzRUnso+UF/X7M3EIrZuGAZdHORdH31VAHwdUN/1P
abx7wCsM1vfISBA+XFSoasEIkQpHt+bDgM3KBT6GlKyFmpvqdqpFGyeprDmz6AX0
+0Nqs4tZRudYR5ohJVIypBWjKimh7wBzWDf7lAUloSIqbiYpYSTeyS/OgIyZ0pP9
QDRsnwKx5cF3e/qvDAzrl3G/Fx5qetJMFVBNDetg8Fo0QVYeARD1IQzme0mSvtM1
C0lV1wCcRlbTGjuQ4n80CsdSkJLqNLn0OkyYWny1ARZRaiFJSWsOwBkjGAClO8rX
lnBpKSid9+PkE9AmmqlGOB9u+fIYCR3Ol3Ny6YYyDCr4VP2Dx+QYz9SP1FKffug8
uZIhluXTf3sKphlfm0lG14KLMEYJIXJ0eNxBi7Oahqs3AiMbvpuRxaRBlzfiTaAk
Fo9HHkauKObDHgAhJnPYtcHLw2/D0BHWiD0l64eFtWI/j41PtFkicrqD0/Qt3Xyg
G14DtMbr0jbeTs6iCvxK0QepBgv66pfH1lVGRWuaw/HiTLBbLgwucK/vPUUSBIqC
/lkRJdKqZPbiTMoSlI/rt4DRDoVOACx23a4iP3pUD8wD/p03bzOPmmbSBPSrT74m
8NMTS64+7V9CPMn0iKluKKvbYf1rZKEU1RwM+xIkf59EcYSVsmBEi9/Cje7EmlYU
29WS4JYb0bSF4pSAMW30rVH4E4YOFTlmIw0N8KFptD6PNdi18PuuJaJJ0kEwsK+/
oH2Ktx0ceDB6IQsM5te/s8pX5xemetMoGFrVINiq2wd/QYjbaF3Sc1qu+/tBm+Qn
rdLDepmIxUaEZsfdtn61aCNr6K0koYFzXMytE5B1lPJ7oqZ1zVzU0zp7PM7frrqZ
/0G3TZx7Hz8o+98sKiHwuTNP68ifTgYh8rsVUreZ+ptl3phdjknRHR5KY/OaJFZc
yBzAvMUxSyCQ1WN+uSCKhTdcfalJldbW0EyKIaABbVizIDOuhplKc6ZrnYHuVHIe
Rnvj7qvmjdLBEMsDtF27NjgF9jVBBFfoXbBNQcscIxcMHhxeX+5kY4UjmVFPP1WG
aZF0qLAAhLEow10rMq++gSvpwgKpwHu5NyQwtE/M6szf/3rQDXOk3hoeOqGS4+Uc
T8dlkz83/BoQUI8lKIj3u9X4PakI5y6ABuUWLLofVEFDTYK3BJPwMmAxkslOB93Z
PXtvS+7DriaNvp4ACmlR0bdquElCSUv2Q+pX8+n1EiS53drdLLSyx2sR8o5GG8AM
DgJNHTHfb/4yK3/n3avQTO49sBRTh51Z1lNwkHlUyEWAkX1iIQQP54V5aQkGXQR8
Biw6h8gntVliwMcfs7SwP5l5zGPifvCaMvdmcRBTALJoGeqEZy7IX3kSzf5HVkg6
qB/5PAKTghmqnGefvgCHW+ZCfu12SyAlj/AiTDsDUUw45HhuQWgNT7E+g2B6DBTv
E5wpvdTKoEpoQWd1vH2pfgSX0Mi+586DmzGwOKmwezSH4V495pGKraeOwPvskoPd
Yk3yBnEOeO018FojOnEF6zaeB1/bM/VZohUvSgU49kNMtEzLPgzuLdN7iybidQDA
zhHWYqrPRV19mXDyUTyW8e74jTJUKVsRydZxpmFzrnrbs6Gz0dZpJYhe5Z/vRffH
FISdKqIpnskHuxPBBMsbqwABwVsNxv0bYhIFM/WMJb0KXXVdmt+0a4JKUpL8keRO
/AwF8mYxHW++N/148vuphGGPksR7qe//ytJm3Yjz/5HOAhvWxFHjUzyjiKAlb9Tw
/EnShbVieLTnAvI6uELvGYf9DQb0o8nUZwtPRIYcnHJMMyGyabfr89ZmieQ7qR9Y
LhJSfWLC9mHN2gEOJ/RwGlJaIjXQiBNRCjc2crK6z0lbDywKMDUwuI/WSwg1GrXZ
xIWMUNBlipIlP7DXMb0SVhVRZeyrRuR0bnVXtuYDJiSPdcUuL0CNF+pZhSBnpS1k
/3E5AUS3qzRQbojKkEWyHBdNHbHDwSl5wGy9KEBXdH1uj+OEmIsXJaB/zfdw7Fvg
0uCySJDLVGTB8f/4xDDTU8wYiynzyacGRmNFJNUIskS/pgF3R03yZrDWYNCvLlEq
H/05+7ZXuJTmMN/MEGz6SeCB9jT6y+ZxR+aTy5wxemTmzG4gOrmfgNdPdnZ4wmWQ
nxR+Li9lg3fC7sQ8LE6lFD1TA+plO2FSI6WhRXp6fhT7LYnU3yIerSU093u+Z5zJ
9HX7YYYo1oXiuUsOHrZNRljX+V14/Y6La5EuGKQpzB4YF2NdxVR1RPxZqbGXc8cI
I4IWYLLfPDRprNUy0Hpl7GkgqUxB7jJJcnHzLM/Kwio74IpCUQUyLnlPla07OhAk
eSd1bAH4GjqEvKFpSx58/hDBfq64+6Rqm6WoBINKCQLGgVEJtIWgFHvnmjZ5x5/g
7mdE6pFaecZkrA0ds/6ZeoV/3o0cPZffGf/6a63AtWgLN/2Vmac15seNrHkMdiEj
iO/g4hDm8NksKpiEVLfrTBm2bCUQeN5cSnBAW+E/yug9TFGnhx31RgW9jxJAgJbY
V5Q25wY+ECO/6A8df18Ptfkx4whQyFt815Bnf23k3EpHdXMcwiMnpTwDPezBNF7v
DzV6vk1VarNkVAtU71cbxbbDLiNxEIcDU3LSM5oVyHzlCZ7wydP1PfbL3/mS/Y+y
aGPPXO78NcdLwMeJVb3CWRqomobYZ9NBA27kQ1XQHSxQfjxvhOatTwV5XGhYLvy4
Hz12xDpy9QvNP8xfF9cJp6oococI5EizgUsz5YWs+YYtWucMM4PmLmXiDEwzncYJ
COW6Cpgsf2kRRE6iRKSYxXqewBELWRDl/RmlgGp0howRmbL9NgicLLAlnxBlD5Qt
55U/eOLNrCHYxNHjzwuaLXXry2/sT2Kfo9Qy3jsy3wheFANKox7m38VWvR/m88//
DxhBzRif40D4dmT5Ch5wtyCtA/KHLuuv0vfzhcg13Kmv8ky7HAqfU6MmeGFnDAeB
+7iXX+SnidbxjUj2KKJ/2s8UPuflW0extVhs7St0PSQCqxetkkLukohxo7EgqcfK
zvXU8CeMMqrlzdTMxe7HNuA/IcZvCUpzOF5QoJA+mjv9vbxNMXTGyq7oVZjsI3hP
4teqaq2FkUjs8rZNnIWWoJqSnMfWNEFbETC0XJeApbyDODGvJX8EbjFNpaybT6Dc
rOrW3MFUu7waQnK0hBZ7ITDa8dXuBvZ0+7wyfXoMzQe/ABT8pImYTHjkfvDeF8ie
o7ScBSk1hB7L0cW3BGY8b6bx/bTuKRul2a+713MKzW5nYtqf3YdphwiSXOJCteyx
1jMNg25oILGq8THFx90zlU1s9nARNt90GLSFIfS/w8bCmkJ1YzcheG87A6pQ0GAy
uDQlEaH1XgY+NwAUpKU9TfQ3bDR85P2rt2BWg0lySY9NxC573UZHMYyhiOhxOcFj
bGOgS+/ITosKKwsNgvQVYoYRYydxomPP2nkzZeyGWVWkhT7itH6KvjXM/sdREZBa
fd4Lv3CzBMTIkxqNRvRsjsHzz3BMlu9HbIRM/Ef3JqFPBZpXsp/nDAQOAYzjjmCw
nTC1OLbp477xxwdX0F3tM64TqkC0OVFh9AXrO1ltCX5c62rBMzhdBxW+SefvYRy2
LFoZybWZb9j5FVQN2BUmA13491fR2Ld+godL3LGSSqJ4JES1r2jLZn7EexZEJadp
RCqDiEsieuJUXzsbde6a28Jy58IZwhmGIcbjRdprBw4qmdIE76lSh4DHApyIKvBz
2E95pLOh3RZt1mFR3rIMnxYdusH0LTHnVFW5bGBE22FPp7q37uHDTNdhXGdOt2xw
FoMmkhQcUSaQADbNK2/B0+DvSR1jmeTJjMOi4JnPO0ebPbkuYGduiCFU2ahmYiC4
k1IzUeqeoZMy83Z4qsRg59hrb+fRbny3X3N+qXAJm4IEOgh6BAkDcIhv1Eo1QfzN
efOw8wwK1F3d/OmxT9vteVjTIZX0uEffem3mrSQbkYOnzpVwf8UefsPDZG4tSBoB
9aekqiJNsPUuVKzKkn+Bef/XYdJLZ2T15KvM0EJ3UDQDkss0Mmr3olqhNZJdj8WM
hcKkgsqLYHuEFWaJUxetq5QAqgW582HDvPUiQVe8EAKCRriGq5O53MEW1foNU6hG
PPPlTsl9ypsy104SdN86P4ZTbRCB0NIj5Q9vS+txwnpX9tPMfpA+QTs+ScPf76Ye
WxPx+nEpLJWp62gSOUz4/8RmyWtIWLag8nDzbF72Pb1C+W8Zuzi92c60hSgcKgfL
BObHzfZGE7Ze6KMaa92anNszBF/XPV2DoQ5pBQc1syYopo4z4TvcXu8VFKtaPsmm
tdl408elP+gaFn5y3iEdkUu/hjs98PHYAp8jFi6h1ZuZPPYq4CUREC2QnHY+04Ij
uLDurc+wBjkvOPW15+qYEIxU0hcrwJaoqqaxHpy7x0e0ndZv5cSmuXD0aWW56B9p
ZXuiBN077phABFC0MhFW8zyBQCPvq8qYa5C7bFrtH8ta8wkoNmRxLmyGIUtUnMRH
ODpDLikPQLhwnfaBhh8Q1+zFKykF/v3zZQML31EXiTN+N2YBcNVxxgH6GcFWubwZ
n3XazRVDJf4uaZ3u8i/FKY36sb3fsaEpeqJaEENvNM8L3SYhm+Go1QiON/15vMfV
vF7TXchjvljTwTSiP79ssmACtH0iJikTw9cRH2gJUn775HGDYt7m875Du56wsWgA
huMtSoFmDJLbsGgYbg0XfMHthGK/rW7+emHpgeYr38m6CttSoxTGhPM0c5OQBIWg
ie1D+r9jIgluSdKvycWh0Ww2wQdVQlaoMVIo2lT4FcWerwTPAMqEOelQuYCxSOCL
SRuTRtJ4rWXxLCVGlNMwmrXDaupeXz4bbfUNqPPCoM1KyOwRiKh4DIPgHIvRekpJ
qT5YzlBabjgrc6T/7AIp4hnFUGKsgkB72reJLeEpIqWYyDdpvbdtI6pYywCmIcNL
e35XCtz6S5hM67/d6+8vWD8jjJO7Jg0a2ME4rFmfS9NOvVQwcu/Ln06X4Zx3HugH
FVA3CrmuJ2MAaxdF2hCR2UL3LpXeheJMGAau1JfcjQ4n8NyM/JBQtvYyNqGW72j2
bM1icIIckJL2A/1oqeuU9mo4ffmnn9C44g4pNB2EGj2vltBlY3kWMBrdBAodKCNH
jide1K55CzFGBRBq71s/AvgP8RhJ8uDWGctVVYsMnH7ohU7HlFrOPX3xeDLDhLel
YK5vr9r6TffC83Aufvehru5Ia3Sv2O+V53ilR4eTtRTBCRPGbZRFSH8LfcpAJl0p
oRf8UeziPFySLVqgT865FVgaM+rpk17lfggtsVEm9rNtm0R9PI07suDrpo6hd6W2
RUmts4FZmn5hCKSfiscuQwRt8CsdWARc7ONPUQjlPcLPD7o75eBISzKHPJKRdZQz
q4e72s87jte/cVjFyqo1mU5S6uFd3rJ+q+d7ZKklhIVxNGqDcTMXgCEy1eSoia0C
MZHL2S7gpF5kaD5+nmGWa/nebmvhlCQBtZgysIvdY2oV02S2nm9Ie636bKiUsVux
RoZkeDtVDxarGnzGFxMYcZer0cJjRTO9PZkp0EWcMavmuSO1EhmHRBCT7v70T/8o
DrW5CojqmB2pZ1IysEIwYeqVUiaAr6StGEpzclwTDFxjBvABNXBDtEMhmnggx3wf
xk8Icz6gYi5vnhpqc3LgEL8ER6cVOxClH5PZG2Nx/mcj2mf0B5gYCmXoj43YpQUx
BHTVpAOs57tGZQe4L1Za7GyCFI78ODtH7wI4Hlh+D5K+IiOXxzPQGduFgO2XjqvR
ZnE47VGpDY+UQiQiTv0xV8j4Ro1EBLK18ssvlAiBmRBmpn9CwNpoHPcJxoNS1sLK
kxfWbRba0lEjA/un+IjSba+4LcgwLTEkJZ9VK7MZZdclv1q6+1uPhXEFKuuTPJgO
IwD/5zgAg/jUEZEARkaudvwvNPxLacccZD+lPjUaKQcbLq4zlHuRsIPgBwtY8NDw
keG+XLCpyraj6vW9eK6ib6NjCVkaUYf48w/hRo4t+Qv475OgvYrOVHwTz7BItX7T
zoxWD3fY/xx/q2PjZaas6TjDMwRBiuByFlLRCkRF46f8DcAwJAVIMumTFJl0ax9c
z62ltoO5ZvU+U6fynyi/L+fmvM8Fzdz+B5R0zHvhzw0EVBpDjGyI3gOl77FNPY5Q
q+2bBVuxkWG1cvwXF4meGimx6Rqg/M1UT5krXicoRpIwNcbkQzPyX2Y/kzz2Pb2n
YY+sA9enH6X963yx82AyokPmQr9/g7WBmqLXTwPfKvvIbHtJiGexbqtP36nge/Tv
8d7Dbt/V/Wfxteo419Uruza5E799YIj/8G8BEeNLXXIn62WCtSo6KvKngGCdlkmk
BfLbpIC4VXbqFhRtLyQtgUQo2QJXFJrKT0Nd0SAHZsT6Y5fjMBzA9gDQfSfnCuEj
AeBdaWzmY0t3+9PDk2cVhMb+FlXMn2eZc4pMhtwU+dgmByulXrm2N3fgGjDxW6Rf
Jn7B1cCzU44jxyqEtmnTM1yvfCnmwCN2CAMmTm+4VlrYrrOpePx3whJQWuymhDiM
Lhrtw8UtJ6aeQqj01VKLzlmAKt2bYmgJb10Da2kVHkR2zgpgACMKhNVaHCtaRSZL
r+KTtxr0W7gMgRxaB4IARteS8Kka6TOjZ2Tq+zwi9MozL6jZeX/vcWSEmg0WOugc
eaOgH+NSvFBOgKKumqzBh3LXDdxCaFdYv33gqHHN6iGZlbOsl9hyHE0D1axktCQk
ko3ga8UodT4wLBitxzWve6djPj/T22UrFT12fLca7UI9QGIGzkCBtISu/0FiUJc1
HaHhdv/vpIHQBm07flHw4esJ1ncjgCUbmWvazP/SXE0PZhX1s/OlKpXuNEtGcB0D
bXG8EwdleZwf05E1yKw9SrRQcHZFca0kbzRR2MAg5920svvk0RQoYF4JnV+f5ZJo
NyYAoOsGAe4fibM+IY69komzesBF6FuKO/GqUEkS2/VKrCgBAT5v8EhK3xRmIgLx
meB7MJKAi9ERcLh47RuBKuZwFuVLSIPLTH4qrCRQyuEivQGLku+SFGRxpArfJza4
GFNlCBqXvA3/WavdbsDKDSgHRNR/TnXy3iPd4nEMh+XoFGC2V6RmjUEyIelnbfm+
8/yfDxhH6xtKVKB1g9DfHzS5o/2z22YtCqbmjiG3dQrDbVrkSzBzR9uqY7CoclDw
tiqUfCM2mW0UiIXnCfnRVlt51tR0ub1Nd4SaYZifrnyQWRpgYlE6/5vXVHubAwdd
OADXBGPhew21qNg1kxDo4vZuN9FTRukxnPYcsO1+7dpNu0FwadX/CJhhqejJZlwQ
yDnE8fjdvaCyltghpTiYOqwEyF/dAK4Eyvt1ESt67wixcJHBGB+zgHXbowIT7JMa
BLl6W8tqbWPl8/xEwd/s0aAyLi0eogSfeTYSN1tBHhVPxeiz+EYoXhWSyc2UdYrh
CuYvH9iQAomvBQgkeHOas9Z1Z68AvSSebE6fi+4X7eg28zXzbKfcvwqvmpGmLQ8J
b5NvlfhSxyihwdJIjuXvnJTvajKksEJ2egK5hR1qYFlTZb+JK11NLi7EoubzTsL/
mgkz8WhRPKB3rsKtWxl3gUz2Tbz/07jn/WImOizgj5VQ9TFoiHKKegnMhixWv9Es
GrSfhHMj80AQlpYQ4uK5IL5fllxjGFZusaWFYySzRL0oKoHQJUKWuWppwwKGgjEW
7hYk4AzzYMeZSKaN5wwgokW6b8MyEQ3v/Jch0dGBs7ttX5SWMXWu+Q3RnhCfkrGQ
SBHM3AcFQtfXst1EpFCsvRATj0K//Ul98JBKjDl2aTdnmtgv0c7lgMuf41uyVnf6
A0foDh7Yx3BxbAVaJe7zgFAMNC0QMOv/qt51r9SjEdzeWk+CYfrZ1bLELDTmEtPb
JuiRdqqIbbYuyJKqoIlyRs45S8TAW6ss1aCrBwu0GeYa1bI+EziR0JIXdW/ULi/Y
2tFB8tXQ0rVF0kacHJvrcq97uK3/xdcVhqQDyAJGC16dxAqvg853j492IZUKNA9P
80sWFbcoy3YLahAXoFIgF8UXly6swqx4Y+6Ieim0dcENjHasp2kPbgpLTnHUawF0
c99FG8Mh/nvm4o0oq37RyonYNGKHPWQ1DSW9p5mggSBey42m035hapcQhtUcxH3g
8YMJteUvtzGftH7EUzsX7soXFvs+Jd6KBmQ503+ozsuZ+RERFrl4MaaUsQtQKdAQ
VBtlO2pLoZJZnQh+kH8FHV4XfpS6nq+b4zYTUG6B8dpgNA+6XmcDjki7cBoMKD7F
11Jm+XnWrcx9wAxt8k8AKAbB0xEPe47AchuI6YHE3JyqRpic4XCz1dOc5a5VNjz/
KTnVdq0ytHDG8o1poFmE2bkxQz9Ju/ziY37zoD8MKORZs+IjWede4QbM0ZyGfy09
idhWOOf7x2YZm7nFqnnWXgxCzlzcYSPS3G6dvs4aXsC3Fwri5cBr/2j3zu779Hei
eKmdFJAm6hxXw3utX1G6/WTOSwZzdV1DcUWaVUKqpbHl1WPGrE6xir6lRGa+duHD
eD/Huy9ykeVvPzvHhwTGxwrMpfmJxehwtwoTXICbSEjiMwqYgpUd+eZ2LY8ucjEU
SzWU9yYcJ/OclpFeDg/EnuHSKHKrzP/ZBuCCQYEcbl38M5M++Nc8Tu4JX7I12Anu
t5HXT4bzYmKUKEvX+4XCucsvJALvyhhGciZAcT8JqiOh1tSHTZDs/EKiEnEdOPGZ
XI5nQZsT+oUR/VA4UlRSGpL+X7wuJZUudvJ5uuwcvcU/ABUaM4JpaUYI11aPkpmf
kriGEkuwFAGXfezlxmIbhcjVsdinkkobzfapA89YXSdPcHERdvCtaOK8sLSX4xWZ
cSjdVa/LQb6Z9JNvE8VAA8i9XMRIMFle4rYU5N//brkYIkA3eBuKsM0+gXz8AR5g
hH9nSeAZVmGAhe3YbEP9fpbREDuT0GDc6P8uarKf99rO0ZvTe404eDXrS9gL7fT5
LiSxqsn7fL7W92OvVsryHIrVwaOoiKxYNHEgWe+HDe37yS+sKOLxyPz44f66LuIo
20qNEGyqHwK068lwsRJ+jqsYB5AzoldCH7havX7mz5L7BXnFeCAk1hyr9aRtBY5L
9sWviQX483wxNWCvkCn6F/RHJu0tv6VzFaVdBqMFXUuGl1VM05LpB9+VR19zqzXQ
la1zbawsCyi5WoTFL4svFT6MNEwpydc/M2xb3iHbfg0Uo6FOrgfXQeGetV90G+m7
2RfBNdNgkPrkF5FmmXkqgM3Un+tOF9FDoWmPTKs6ehJkWT4E/JGYS7emc7r4WCIX
m/9lT6iZbMHKDvxrEz/VQYmId5z9zv+z6f9HfncLab79DIALxRukOnXLltAX2kVL
65fT5kbszRFHfMP/doTbQDU+vYOGnvdicYEOo/ntHh9SbBj/jMFidnGUKRaiCFOx
7uoCQDYLakHZpSxM6RZ9iMSHJ/Y5pravHkVbsgaJLuwGxXAQHnYRX97ufLXoT4Mi
mGtl9vrD9dPaHhiK8QF+WaJH5V3I/ITQKTmHalHZ4xoizB4lOEkBykr9U1lHRu1M
FELVrtMJc0zIneADR5h+rTXHggbSg6WpkGjQfv1+4+xe43iKydelxGwpn89EIRUh
8HBLF/aNRwSlWN7G8MxBpclxQJtjY7qKqiBrTmWD8T2OyOPT/BLXouFbnp4kjHjU
yWvih05DsMXbLjAyodKrfublwMlFa65i3rMVHELO5l8RioDQFsV4G4+t0+nDTR46
hvd4jtWUcfJbUlekXSS3QWF9zh0BEDgdm/z1229iArHI3ztgdIzxW0nbfaFXrw1D
2ikaKb26JHfq8jRlgGPQ++ILX+SMHqx51bAXUu6+E4/WfKZHk/ScQaFK28J3RC6R
/CM1wobmB2yjd2PlPZfKcdOtnxELoZVdfZCFe33dsK3hN6sKnzQKNid/oMblewoL
sk4jx+ipjU2DBsaO+S+mfhw3/rJmMCqeDXOa1bhHv6nfqtrZQzvt8uI7ushViYCc
xsmcVkEL5imMLzRQjdp51caGWHtQV+ljwIdSJllwafDBhMKE1AXkJiaAiSATfkF/
2IZ86YO6+2MbsChPgbUcGLIGmtEA+UkZ0UgXjf4LDgoLoZBmIE4ceOTnEJmQqJft
2+AF2RedunBI4unXbYZthdirmev2BoV+B9+ddCvC21/yYndN6E2sLLImHqQLb3BQ
bythpQWVYucLDaoAh84WPa+8tJnDffN3o9S0XJrUVydH80xPOOF5wlwEDqW1AxYJ
x17TVuXSdj+lf9J5gm3x/aDg5wDfW5b0gUPe0AE8LaSiv5dquK0FNz+esOI8oMkW
LnhhJz8Q9dyJtMPhVlff8VZxmh6TD5BlUIDv0qlSIP1vbp5fG8ORecg8kfmrpXmy
bfnV/9vQ4iT92ZWIPOQHgCLgs/RJ7YF4z2tjs+D/RzJB4D0S85vgXJxUxh66ItQe
tRwHIIT56uG4J7LO/MdQWmXAqgY+kkVirLnY3DsurN+Op7IRUhR7aLG8jDKg+Cdb
+cZygcKZwS4ZVF80vgCe4XH5diNHOPFAO95rnzASkFjJ2Z9ckUyLz+Bx7U4VUIX0
N+2lUREdCKK4FSEai1wmYpWVymnBYLDRV7WUekW4hFanaedSU1u1WhGRJD46CNj8
KzSvpGMP9Sv+El9vxQKa3/CKSzBrchx8m4U9G5Dq8qZuEUkzGLT5afv7sLdjmGcH
wtyVoldp9rwZlXCOQFRceG2Vz39zUgSoEMekdCj6/9M9qoZEAki8eFGZKUkdTcTM
OINc+voCtvq4CfNlOYf+HJnyIHmHP6dSiBDzBfdUZ/5SXScWAliIwEjzhPZZghco
xGCrMMd4WooIedARxnTwGn6Hjxo1W62CKBIR0oGD7GemZqpRsElnslKk5K8+4LhQ
dAHx87Lle64/ovVqtpKORpdw0ljTZUE2MEr5m7SilZjOR7EO8wEDV+/5ymQOutBy
PrPSLpAq7/k5vfvyOwwNakFNcQGypiWXtr5MDrar1Gf17NlYTXrzxG04ozJEWlgn
dr9jt3y4T9SmIz6pfoCJ35pn95aG0VWLDQ2LD51O6tMK0oGb+VSiDC+Cf76GPFDA
1K5f7eEMmjG1teiRV67ONjZQFi5T5fO9At8jr7PWlrrtM//RX3S0ypIe1xlPBZs1
sUdRHWDDTYS9pDV+dCkM14MsoDnQoeK5e216amqM162X8S2MNRGjBWy7lQ+w0NT5
VYBDdSauC3MQQ786y73ZII6YQ9RL6+HXZo6g2SWUdxvEYqZMA1mDi5Y3JyfrFMYN
mX7UbctVMOWkaOKPFNYaPGba2D1bPMv3Yzcmssg92MEHPNKKe3hZzE3wKNi+X2G7
Z7BNe3m6/jcxXS5FsokTGm3GK4CUaZ8y3DplRDJeNREryur84hvJ71b0Av28qhhq
8N9Qz5RmEFijFlhmUrnwDjP4CUfAZRWLO4bap2q1OSZ2rzx5or9XdWWwVFxcLcWf
2QBpfgWXr8Xxv6WYSxoBZCyKiex3x1g3ftwBNKppSuR1vwAyclVwLhOq++3jiUQX
MzMgWkpOmBgmswJq/8X935SyEvB425wITG7luNq8Ssv1OC0KjgRG3nH4CQ77Xuqy
BPpHLK7kh8FnXTiRwZksMtFmsdrv2CjsElJxlaaNlO9VZczkP2CyWYO4aXCrzbpd
p2VQkyNHeqt/+gTftnt4jRcHN2UdqbytCL1NxswEGXZah7IWvjTYZplijYAlTqBP
zm5I1fVyCxUJBqhDTmpnE0lJn8SVcAWI5XJavZe/n47iFM/zd6NLdeExXHzD3ur4
VwHAwARpy40t8JMvk7wvujiSO+lAlg5Ka0ETh/aTXtSwYiO6DIhpT5R4E8J+niFl
NNr41UjwSElnqxReTAxslor4lkyKgq2A9j+uEncfM4doZjAw6Vpg3xA/p+bmrC5S
VCNKWPfsJ9VqKoV8QFhArxQVy1kxGj/bNYH0b1SaVqr8J3iUcRiGgkFNmhOPepfO
75gl0H+oz59LV5qO73hBzvsYC13TCUXNhUSpQPMLAzf4m/iFYLD1/ur3J7c5jEkk
Jzx4DHOgrsNZo2pNlNfZppjwWyTZy9L0EZQmQnttkIhVmLiNn2f4Gewq4tTsiyAE
BjBNawJrct+ucxBzw+lSvN78d+ttp3+bfj1YrkeGbAmmAXWL8mFVAePsTicHw0pu
ANZ02yGYtZ3Ay6QjGhiKOPHNV2y4x/QmenaAbFBsijeos5/g78WuOIQY0ahhX1Qy
MAoSu6bhAOqk6NdiSfiwg2FawykM4QjHygWkN9gfZ/N20IBtkjmZtLKHbwSFLeFV
GrYFPlKFE2c/id5HF6LO/bc8E2ZgkY3S0y2uwVBfRnWxUG3hAnG9nxQQhGOiZtvm
2yc1GrND8uRA4OVFRCj2PoxMZ2FLn4nYdOfbNOcCn9+zdAM26Pl6kPUInHX9zz9e
lpbAGkWnDD+QVCI6BE49nHXYDDmA8m7E8QqVGZO9d76UB0/Zr3yFNQn4smTvXS5I
Dn76HU6zKHtgG4WIxnAJOYlcZSQh3ZL2WCPxTzxAfWjYRvdwJkFta8xIdOyqDucK
KnOIRB7VYoKLDeHae/Q2dNn8ziPl2wFwJaf9fRo70J5CuC9NfL57BFnBLCLKbsRc
KKBpoDaO2u2RBBlbcDNweXgoyH4tXALv2eli4PH85lfcQv75JXrK/d5CKr5UFREZ
DhchWcdIV4Hu51iscQviIA1HHYjPjoIZy/b9lUKNJfda4+Kjc+PorgrnV5djCnOJ
TApMXt4DltwvbJ0mCB2FqgFXY7RK+EbnDqPcpXiKMpZSQKaoQAtY0mze8EBNuYuB
T/+i08roKQXWvUtEpL46bztFOs5Wf7GAXt6YFvbeDxoyUizLXewoavP48o7D22Zn
C1vvzjsQxvtfLNbGTIys6p68TsFWt7PQDrENTSrjzJJqmx4Yhm49NQwsnuetgixE
RbsxinGMi1vn37Pm7oeDvxN8oH6ko0MMjoYCe2cw5rHCr9FtyiU1txceBIcvKtq0
aFzjO1WIrdZrdrHPSUgo4DAVwWpd4cr5QciSj2a9IvSQNUuARTfSqL5Ut/NjYZiu
xZZACg7bgvliKFWn6NvestrlB5FxG/jU9sxVJ+mXB3jOQzzVJNFop4CsFeMnfbmq
2Zoq3jBQT4fgWdIi2QAIa8/eVKGY7KZ/hPrZurQXet33VEB/c5Ynhe3aJloeannc
hG5cfaYH/wRPMoEL32fEcNptIDPTrBMVes7cOzokMeniI4ZKKePVKK3Uhx3aAtzr
uwtp4RiwEA5IS2K68uyvUKHhfGP5wnnUTqpuabyAo00VbZAoVcg7CmXqvLqzwbAl
E6Wg3Y/+n+WYEtzkIjD5PProBlLex6URdfA9L0oCeuF5tkBYl6JQYi6ZQ1PgoTxA
54iH4XjDTa8rL4RoZ0mweXKHKFG/VO88M1Fc987Pkg1noVWfRlbXCY4IxoOSHo6V
8qTnSIxMoTgIuIfFXz44d78PeHTdiPyumuaZKu5F/rSBisxZZwT2dW1deGmssYaa
flL7lBD5SlfcJwe6ZCYjMC/SRKD2+2qJ5It3im+Em86D0/02Dn/V1JtH/zuPeRD1
Ow5eD5UD+0oOhAW9ZCViYPjDe7Kj8MAFeRASq7jbKwRCB8Ty/oZQGKNe4rJjjX0D
14+3RpHVPsH0RjsV/O4t6kJLKfrgJ8k7RM7NElEkg1x+dgQ3Ox6m64i/qsT4b0i7
EiFycNgRxTC3VLqr7cqsTQhfykgLoBcX3SAhpjALjpeaO6vwIuD358JtOBgseem7
QGQhoU3U87sPCIOYAG3c6Ayo7ZIChDC4nq1pl0V8t44hzqgMh+fr1wf5LxZCiEH5
IHu9FCFmxDS4agoXPwvCAOLMa0KLejUYNXLBOvCGuCSbPEMB8AQOnd2cRRa6sUmH
LtKDbmwbionPGWd9zuYpavxhrAjWHqD9mbHxeeJT7AI8mgSKny7EsA2mOCYrMH93
OCWcnsyaXE2VtBjDf3hDxx0YFet0HmfpCmfPJJ7mkL0SsDwUvAdmghJZ9HCdLBoo
rtJkYdmj1Fdcvv2XhqkJZhNcuH/VHiuBtYI/R0dEYciW3xzmD8iOzT7h0eOW8kOt
sGWJgzrXSDmWMd01BO94u3Fu4j7qUQtID+aBTywIA5P+MZJrQhnceUmbaRX3JhAV
/HU16zFwU0MYcq4G/6zLE8PrsGxiId3JB0olTiJBPVK2AWzyTdwe9+/kd8HljGyG
TtSLs+4VIFuEDX7y1NWhv2rqIzhChSjkBC1dvJz5SZIHI6o6q69C8Q6Bs+rBU81l
zjPBAsS0WAu2hcjpxCQnFFj6zhSnGIbTRhGsuvFnV1wTgenFnjJhVnxvHiGv+m49
epLhvVjn2M9RDbDAZudZKPcJZ2aPs3U+HV/gb/8UgN1dtOM+VbBGkpABzFxdxk+R
m4DZVqFJpFeHXZKADLYlVXxbjppTDnC4F7/BSjUgffwxMzs10kemKXSuqfpB0SBa
XDD5cHXPF0pWLj/LAIDlRvJiPKJ1l5Ma8+mVRenrxwTvtMLHxWWkh4gqdUQGaRno
ueq7KUq6L5UZHABWU1j24jKT4g0vzzCJ7z8zdayWMEkfTvBlPqpK+KFZ/pYK7u1B
lPXsWOOfkZA5SkP9YAqMmEOmC1dQkn9UadqORMNHrBlmm9y0quorIxm1filQ7BMI
kRdJzxBYi4SFZfyGwxGRDRxoEaP5wdr9UojyIwp+xgNh4VWZk7Cv2dx59LXNwHmu
bLJDst02LV1nCw/H/xwc8yDut7FCw4XYfUr+/236f5bO0WyKtVFOnv8+Oa8Z1ZNX
PmQMEsEePSmOxiuJnGcwlbSpHWgfHMxHY5W8pTfFIolSxWnPc6yczI4mttBUiShZ
JOpPpDQnvsEFX1Ft5KZSr61Kh3uFhepS1F3QsMaflQfYSHupmN7B/MQMmVJb9RGf
50C5RocJpR0AJUTyrfUNAlUmelPkgoWHOfSOqZsyZkVgmJCbrCs8SrPFlZaVrNg6
Mxm8RhuQZ9aeHBFi5r/p9aOrtXN6cjCmrZSPd0+C6HZ+dGDRFtV3H6WYcrcSiN61
YibJkYydKK4xWjOLeasHGtjag9L7g1VVTNyxMW7kAmIOI5xjppgz//PbC/LuZ66G
jM6nd0KLIsvDRIG0VUkg5+G9lKct3p1nFqTOGjOgul7zXjDJsFRXPpwp5L9azfn5
QX4tl45AET8YUCgKD4dLy0TaS4oXCerVMlDfzzY0hialtqT9falmKMHOXkboWOSJ
iATdcG0D4okK3Ck+NcbiUR8CpPtF7r8WlB/ddUYviZDOwdRp6JlUwN/Omc0PaYPN
Xruh0Et/CtspX+ff89CK8qH414MuL+s58gmKImfgJY4Y7O4UY111a1ECh6Y2z4uN
N0GHFagwBdJE2rrff4xt1jtlKXOp7ov+xxbkUhfZiElQsNsLhPAn1MuoLwZgso4m
byQql97FZRcYaiPOVzRr0aFPE7xEjtRbp0wDqmtibF3K5Fd3Wn4pxRHHN2BJnFp6
OZzHzHgyJBOaYyCQcSgRvWS7MzUpJzHHBvIoroPD2/7EdRzdOvB8xrpPmTz4R1Zw
/p37rW0BkfoUtE/SAbh3PUDAdzts1RbFS/l6rUUacOXbI+QzV4zKpyfngFx9Cze3
G2IpDkCGMrP51Tbir3GdB5K9Vz9mJiC+EsHt/mZcxDZwIr7EU1Te3iIYThXl8sdc
/0P9eV1VXMtL/jvYE20vIwO0uAAsv1CNrCTNUU/++hIwziChaQbKSOZlklCh081/
Be6BSVa2GACphHxhVpYz4xtIC2ipOwyRR5m6Bk66/zbysaT3TRpAE6PVG1Y+v+hD
EKDrb76nbfuwLCNgWjourJ9UAAOIZVQNY8xEv3ndkbbrgUBFUAc5wk7YgLBqjXrS
zO7Mn75Jj1ZXgZRFs73XiExyGo/KhONNLy2p3wa2NqV6cguGEmKKldjfh1Elr42d
HdqVZRDbXKT9WMxhSX+6PdL8LWpe19NHwRzOY4SNknAx2XXV9x3VqdczzBveIvZ2
iU1kzBBC9N4ULRGDw92Rc159ffAZ5VRiHYsJZmvKQr9l1zKjE9yUKGG8xoNsuMQL
/Om/9NUrVBwpGC6VusSTBATUXuhf2+J8F1JJIllaPMVsvx0Y/Frp3Tj7f06L3UdR
I71/57UeIWcOMlrZzAnk9vYbC6A2UyaWAMkZI2aCZzuEJmKLICNlouaRAvXugL7J
HsdG6LsbqRNColCSm8fo3pgiSw4SbgGhNEIJgSe1GGZhE/b/8GqMW+XUa713zKHt
mDP1K0cu+EcfYOO1jrjsA6L486efglITscm9/PTrSWUUwlqZUIRhGs9EiNubVJDb
Kg0cwBheNfkdrdLskpXmA9Ee93GDp65xwgZ0Rs7OW6mAp8AqPGTnwOO0KMTnwezj
y64pqINkKVbgiRcECXz2CXAfzDpLDbAVcTKmQgjdwy9NU/dUBdHjQb8kQH97XK9G
xgDLIcPMEMB98G/nvh3hDuU+Zkf85rtnz/rzd8iXme0LXrpflWO3cqG3luGbphcL
YZDVAtCiBN1VUvvv1bFaA3w9glmf6UAFQdXrjJFAEpufGKLypi7krxAV1Du+BOYb
I3WEFE09KQAt5Ak+Q4DAXSnhSb3P2Xw9e+feroh2ZUpK5wzZVpW6nEksbOfcEi/C
Oyaoue3UgtWjaTwBcpnYyBg0k7KNVPZbdT0WhyLDSp7tgvYvx020bZcsWhBLWe+8
4GTs90+AFKDfx17yZvMl8gXN2/4y7yyZps1haQ1dr3r62rlo0khe2xaGcb4NLr4S
TQ/v/wU9n9ygPvsHoJXtyeUdHkyZ9PAufzkzIA6yt/0M3iFlnteN6IHkJUeLuvY7
T5gxmONU84jIsj9i8UsYW2FnStfhGzk3Z0KPW5TkDIQDiyK4GVle5dDkJWCt6vts
4BRHorNJOFXSgcIP3QdPKmIfbOoI4eRps9yM40YW/Uxmc0mZtxnGWptPt21UOZbb
CNCM/XKrKFNJctUkG9cRq3OCfF8vgx4UlJmp3Xiqx2Kl/L9g/BPjGZPIR3fTfLfl
W5E8HeZV637H/doqIbHPSKTIYvdVEXJxC89it7G2JTvzGZwbADOyue5aRtF9CwXa
53Fi8sY8O4bxMaNFQGeVzLVlf6qMTiDyAdhicJx9mKU3Fy4Li9X97CQIXRVQUhVf
gr+2ZzPqTzeQT0ttgxGqYX3xkWlPoscZ6h+PlCz2mRXbmbuSsg9KlOVTIJ80FjAl
VqLR9/3t6SU1W8oxCwBBLt5+0Ghu9xpu9PfCacZAqyxAX5dIkVjbbbXwdOmQ/Ze3
ioXYaJ5o/wUhBD2pg84sPAabc6cUxHy92a5gN+uSc0SZX0lauxTxb1naI4FuFeBD
VK32X6pzVMcyGhfotKikcdk8SKGq1+kqsZXpfdgibP3W0HQUvF70Ea49MfHRhCTV
WiwPsChD09p83EOUkigCXQZdBwWaddyrjmnYayi92wRy20GUm8uiHg63A+Du4F4l
/zB5ZPh8DzVNjKtZn2oiP2GL9qLPwCNX+qZW3kTWJd7HwMl2KbYqfqdyV+9Bn/Sr
DDNQUFtiYDNNcogohi3g1hi1nrm2LZyG8o0CsGViinPEKfj40MkLjUUGbFOQoZAt
4Im6ji0XzMnFHilcztu5HTxNRnUsH+NI8dGbCGPMK2DBY/3EXQpCOJ/hLakZ9fhS
udyAX2Eaw0tmnrC/geGzwbPkTWHcduIdH+rUN9NPfALGxElgWdlp+Yh/xugmLX/y
O3el9Nynw/GKhAH8k7BjZEP3c18YfXWxKPgeaipqTlV9+Qk6nR/Yxo2nhbLJubI6
1BFcFa8nI6Me/1VQUGDeg4ohHRM9flCvD0Jg9/WQe9faKZUE1cxtSmBgDldg+GRQ
HAfCNjiKeucgNrYBWVYt39jHaEAoiNk6D9toOPVOGPZ5HJiMXVV9YL0PbYoXWfEV
3RMftxOOuNVUorFXHcJSxeJJrV+NeBVp8FjcVK54NPNqBA8EJ2r3QOUnd6tsujEd
i/IAIh3AxvpU3KyB9R8Ky3HDGSIM+lKM7wvv/Z0TK5URIFoNbCsIllR3PAWszo9G
79jLhS3po7DaBxX6mHxnGwZslq3chvT5tdJOwgPcpiUUUEKQdRX41Dk0bX3Lxjvn
OTyaf+HUmUhXoADHaG/XgFykZV+e/G/zO1gdDl2iREqZ9UdqhboOSzoJOkO52uL6
kYb77TdHGyNBtclsbOnekhNG9V8vkCSBmTAHqCuGvNyJ+/PqOhhzXhoFsoGryLVm
CbGd54l7Dcsa0ILhOYjcLke8d2pgegFDA/xWoOwSuYpoURBwuf0RdU2u5mmBr1Ck
U1krXKoAf3rmRdxeYrLrYUNt8NWURW34KqqkV6JDeVSIiFaVYlDl6+PbPpUvYugW
ityWvDfbLrmMC4pQPDAHwhRp2zrpFd4DOxkMgjvBZH+qfBqvqivAS2ZpEuCliJth
lEJd2J4JOLs7v/6SBVUs/DlQI7JKQDho/JYB0hhH4KiALTxynbQQV6sBqg3Gsj3b
MzZMHyTGbhUJ3oZmFyDss3+QBF+TW3RxhQYrTHh8D+oUCct1HjZyKWYhFm6iIYWI
Hv0BEB9RRSTQpjNjY+m8wBdhc5mtE1J4gWmwYaai4MHPkctnUH71TaI418xMXVIk
KET0ePJwEaG5OCpLgssRJIM5ijVbFLu0WRarkz99Hkcio0V8Z/0j+WdLpTYyiIPE
jCHuLpFbYBud5vZSRIqT6bKNnVQpSk0Q3hdFuZYyzCr5JfZB8ADsd290DoXyzRQ9
oeiXs+D/Afy4K/H/XVDX37fm54T690oM9S0qfxgr31I/hA0FBC4+QjLddBIZYnMO
FK00ZyotAtszn3G/EhoM7cFPgOkD7DAICVn26/kItaTre74Jf9jWOFQQ3AfnlkpY
ljoaZSSs/cUt1aizkzw3mpvqBLNtXCl9Qu7tvDwOnIFSNyxvq/u6n14383JmmPSw
6C5TuzmA3xeXJ2OPFlVcCVVU0ZkBMcbq/WXnpHJGvTL0VJAjIaJuVZmsQpUvrvXT
KPV3859tUQVjDgnJpPXhyMiD+VvsFzfaahuy8mIuE79iUwB5S4e33KG3z10NykiE
HVdHCfLm9Zsq34jNjjBpCmx4XAuHj/2VvYrSufZ6/axQ1y8JXSwAsQPFHfoaMgTY
YZesLJqRdtrnrTSSEN1NEpTD4Or5VxMZ2+akjHabr6xF4Mhi84Kx8FkBYtBhqO8A
SeuYkKe0ZV33Ww8CuEHtmesQvNJ6oKLhn690HViu+DKGA5Q22iOeDS2x3dDezZaQ
fl7I0I9HlUeCq97J+3Ib4ds4dv/wHp8+0IVLRL2SHnCJZxVIDmeDGULAmJGW6TRa
F4y7V5I+TBiAGTBGn9xyI7JG3FY/frMr37yFvAKvBDOujDeRSdI/yA+0afuCUZS3
ITvWZ79glOxeTNJPQ4qUsOGloXySEHlv301Di5IA+buybV8HuSXMOu+fl+22g2sc
7486Q0PbtiuSJI1ebY7ilSQPRsmIhw74CyPfaPZbXtZ7R1ZiR1e4G4AFfffNWeks
1s0o4yRjUxw1PAlmRNkqMgid+KLCUAv1RLiD6yHwQWu35iVMSxfeWtYywRd/cRrU
j2Pa7QaS/xFWY+yxPRBv1RgufQCXhWknygxadB+rvkzPeE3/ZH7fZjdsbgKryPZB
4UclHR2++jozOIpPz2zckKBF9a6VmbumjiNMPhn35xmtqPoBBfHUqkJwY0V5xJ3L
A8fnZCQIsuWj9rU1HpZ2wjnfqmlEeYCng7BNfFKAAr+MC3WogICxtBCJTs5NSVYU
NMLShBCG+p4J5qHWIjUgV81H/oR27UZieuejaQhPuMxkY9STIV912RF/wnaPc8jr
5kIPT+s/9N/jgU+6AOw+cKr5MXSSge5FUzZfRUKkIODq/feOAJyzLH7hKLGgdQuf
IesIgeXAKfMzq11yPhpc/pA6YotwMT+mrW0WXK0+z58zdx+s4yDq1H4aVWuq9imO
g2cxj1B8VTtIvPoBgcbyLxIaZJVKNS4Ou0oF6CUok+GXPPGXqvJcDTYmmv6LbJAC
bHU7Hu8Jcwt2S67f9mORJkMilSM/pZ2cLhnLfkv2GCidm3xYiO+GEVZarXo+/G4Y
RU+neRaoqzdaiR6uRKJC9ZiSaceWHHURfVFfp7SCj2qRtKx1GInpJyM3TzbDg+Ei
aWMcGWVd4PyrfRhOZg9J17eKoMgM19zovj1f612CagsKlzuAS5oHaL40YsIT7Bth
seWywSxWv9/EECqlflMLV0vMjqTQjNpvxI+dO3lgr33fgp7Vfhx0MXKiuPyR55qv
Vt22wuSa8jlhjE4E5iHtMI0EfrGCjdM9bzJs7RTe1GN/AGNAZV5aGNByhe3Z5q9Y
lhlGQerLjLxLIM7AEGXWIOnq4KudUSw2N1cDPZpJENytMXuaWohaeeIcoAjSjhJu
/9C4xRwtYXeryjT0Kn8lBiPC9KY64W9+bEdE1VBqilRn1vwe3V7Jn6FakMkM9Pv9
ZGtMwqevuVV11818XI+II+9chwi6Bhuuzu/8nXEUBODiGAI7epckC2fYeXpS4c7q
Ne+lsi2kr/Le0zbf/tqx+IO3J9HJxX8lt68CWZS3I54M0ABt2v45o2YNsr+/Hcul
Z42po3w61MACFcsbzPr3Q1NeI8RzKgZaOGk8l4GTLc0lLc4HC0ySNSgm+aMan9Cl
IwuCvl0b4i4Y2vOseOrpMkmFsHD72ut0us+eSzyX5aNWaY4nzsgTfN+DMXgt5OKu
meCVexvyNPkRa+Qr3qp87bKewVgIQQUWjokcQqoAQ5Pp8jC9xv62xq+3Fdpd0RZi
FKrCWeNMOmtfJNZ5lDSLPwm9uTCKGWGnIhJdSnYVxmr9JqSb7v9R8qcENhLY6z6T
WriEqPUC3i8Ff6mShy9HPCvefff/TPAVflNPeVHUJSLiyIrc/pU5k5qUf+TysmAl
tEcCFE5oJh5uQq+pDCfpuhuDBIYpQrX8FoTXAsmZXf+U61VJceMuldXHHZ9ilEfR
66/n5XiOQi+58Cw9B/8C2NZJnWN0kqA5IdLHIHER62reh1Ot9yJKWqpPCV9V9+8w
MD4cpe+cim9rfCERO1IqdAAlJaQx++5BjzVZYDYszBxfCELs3x4eEwvRnG1ft5Jk
tDTNNtLvIWoyUigx0CKq5EVWwWUQvbTz2BPQuECDWZd88dBilr449blT3dzmSNSB
fIa9BgcfVCQhozToYwtcwGwhSLSTyFBdWX+bYHSQJShVmB/sU+HltU9dy7268tyM
AmalkuXTSVQjxAVKZ2Q4YL5mkvbE1+P7kHR3CVY3XWuLJIoggG4OYRDSONKEBojF
e7/R/t6k63LeliGsDEZ/NOFYJ+wQLRjrcpbrMPtdwtjUuZ3MppHI+GFLt4k1iDa8
Y3AnSciMVblhrAYbZ4c0bBe/Ool9dh1V0Z+iDdONbJwVy31S/so2/MD1UQG86bUv
erWJQUQMKStUyoLYH9sb9LtYAAUTbCAw8UwMWwGezypmuvTmZrCe8ujmojLkb/UR
ojfreb93RxYakuPrDqRxHcuJcAArXKa11yLu2e3HvfxGSFuieWJhJPaP3wTtaYlZ
q1zJUjFKsknRE+P7cnbCWRp8FUG9IDLKsqix1biIKhVtKKP0LUBgIkSb45+3mkzp
6/9eplnyg7RyhznyBUGFqmoDmSMbN+vmMxjtYGbz7RYpAFwanM5lEdGC/zr7t043
bBhX8BaGfV9EgipajKvd0E3AaIQkcOWrqCsvOTb7IU9gbj4YR6yCf8wfEtzgHALC
1EFWm4q+rSziz3PvGgO6hi6MZxMiRxpOM/yFWDZZlz46OVJBrRPtK9CClMil0mE5
/zsZ9NuutO50gMAsl5qfYlW8IfSAW4Md9u18faMe1scPHuZp9t/YyoieF5B2XQ+g
ApyM6bVvsWxJcMfSyYkXodUs4Yv8H2zn1QplhFIrgWAT8oSAtKZyAVzUgZgz8qbT
qINHGeRTyHv3plbPNw25N5L4c2ymjs8zsqgoikX/fCtrzopH6Y7YMo1XRacku9xk
Ml3sHZi92WSCV4ZNbQXJsSEngy+YSCf2aGINtIhejCvx6xHplPfiUnvEwTKUvNCC
3MlZZXq9+Dn4MBluCs1coIxZqH20ga4Ex8YiLv4dt4O0PiQsUYtkmMzjnjZ+sFx4
o7J3ZzGJxaRLT1kec3gs+Dpl3crEs8VVY4A/ESRxZYbF3lKw2xCJZHsSgz626jkw
HQOVmzifnmf8FT7q9f69oZxteGwtZbBEod/gpd6qnBzfVX/79d85sTVPnhKuyl0I
1df7cdhVomblPPAaEfkTr8L2i8yyn5OmZxYZyxtP0/KfggbKiUJsTB6Ynyo51Zbt
jspNpNAK/wk1X48A7nz9g2UtAnwLDHqLA1d5JwygIcZhyzW0EzR3X/180U7qJ+ZE
y1pPITpQNWDxnc+eIfudC2UitaxpJhKkuSu5ZeAMEtzBemosFLhmtUmozgPCey+T
KqISe7q1PApXDDoqrp7KE/sCEn5Z/6cLCFpD/wiBnJKBvvINOxDaQBI3FubUOTxg
a5oS6zGUNoU8igwkJcRV2eajRqt6P92nU7e5E9KO7yR26dLzfM1TAE+fJzMfAZOf
JF2p5Eyvc1WPyEhwfYEHQl9gsw8/p66cKQizKthblaks5biEq2oZMHrt/jDjguYy
yW1WKWzXVIgXVAcPDCb2aL8y3HqIIAaB2MFdojqgJJUUhZgQEEp0Z9hz+twqcpFM
QNhg1NwE6YAVCXPYVz3wjM5Etw6kFFd4+NovSFLNUz4HU7ar3G1LHpASLySsdKdU
S+YoYXxZq0awY5HzBhFLD5LEFfn9oUGidu6t9s1EZlzHQnnWgD0r0ionXy+7IpaP
9G+AWmaE5rRB5l1EdVASWfiqN+e7Tdtz5OJ95DwaL0r9ZJAe6/gAoMehx4EN0rwZ
9xkn/N0XbdHR1bsvjIhZYxwrf/o+7eGNwCyb4spDCOp21k7LpF3t0GewHQKhEqSI
7szQHYnBvra523ck8YInOBAbArHfSzjs7vSBAaZxVoJ7+beT8J1Et6vgQYPkVndd
+IrOAM3liczvqNt6lfO4EKk46D0Am8ylN9zKj55WJUq/8j38DXPVeHA6N7M892+u
lpPBf2EQd+L2o3bxs/JQ424lSz5DakghXECnJHcIGl1PaujcwPko1zos9/Fh0xFZ
Vqn21j+JlzqAublBE87pSRQhYQ9gX+ylbijyX8URmhCq/5ZBw8VeH3dESXIJY7Zn
j+zCisvaIVYr8uXtcL/7FMb7xYu7tjDAR7mYJZ/tIIdczK8ryd2S8awIp1qBJy4E
6Dbe2svpzT4c2dUBYY7SKPuTVFfyOyLkL/73beZSnJAzTz82UHIl5rm7uoScFT6Q
3bLQl+TYvXrbSr+OPmKdMKs+87igEsrT/g2u5hU/LKvv0WI06d8eY5hxYvS/6w+e
pI9f8rBoBl7VcgdV4QF74SQAa3pLCYkDiVS9+6Ip2sR4KxefoqyBHmkwbU48hXhR
LeZdBmH3bf+wKTlx8TgH2n74qdNHuVjXhRB6/FimO7CVbsPXRGljf/gRxDhQEJiX
uNi39mZ8J6r4loQ/lkSWDxdqBFKlDO7zAnujLkoinS8VJsji00l46iKR3Cps4Gsr
b2CQGJVci+Pck43+kVhsxrEM4ed5f1FyK3nWuG6TbXWP5uAmodSakaneFFZ1WIGR
s3TF9FxK8Q14xyWCJAb9RJkKaw0hDMAWrY0OfMcoSNzJPGf6iG6+cR/9rwpQYYhF
PzGu/kP+sJGQCG5A743Z2xJfNfkMQL0F8zzy3xt80j7haepGX0Yk0sQl9r/TnNyC
5G3JrnKnnIHl2ISjmSP3VoOquDCnMrz7Q5S93QfhjESeWK76nxV/CInkU/nNX6nl
Be6CdGopZOUAgycTw07YQYV6+hNul9dt12qs7hOaISmMXddKvIGejM2YnyxQ2VJl
lt1lo4lbILtaWX1SOgo7DcrekeC0lmaKwtPx3MoSaMKGASCA73c8OHUZbhuvJgIl
fAskJhpdePi9/pVGJ3IQVDHMv5khF2rzlVAY80f4ruETTLEf9JYWkFsbssUW8nJv
C5Nbmvgbmk17R/phIQGPiESC0B+bI2NOjivhkRKsMSK6tXSd10gqJH7Gfz2/TIIW
6g91/tux+sxeBS5vBas+o063OBSO/pCulmmOcjdHzKcLXMN4a5sOnTEfmEh+usTR
6xwCf08JPJW73LSbGIb0eJ1lJzxy94HNaLsj6zH4TaFU0FyM4p8iVCBOYmQi2nPW
pwq7VrfjcI4C3qZGizxIafKvS8D17euGoTYORRHtaLQbwN6oPr8qytTwEgdqFmg8
/flA9hUbadYMdS20jZHy/Htf8LkFQ1TKLOm632TTRbSSWpYFvUTGasERgKrY+725
xxaWhGHNrucYifaKanQCyTbtFxuMxtrI1Es9EKYUWZZiXvclPltIJdgpn4lrGiyq
bZIg83F3EHhyY88Lyf2txColagGmWCE19oDbj4a7H2N8GW99/g0qBCA68VacP6tA
qcm0ySqqQvnumDtC75+tel38ru3tGFjlA8psUdxMNBUYGuc6rs8/Yo2+RDtWo0qW
TQTMWU7R91D6D/5rwvPgVP2hiKT9+SVo1mhHU7V/FfiVBFApe/ajGhdSqCmbpzGc
vsR4KlHvGfh/zlovWXeZDoMktSV4kgT9YyYIrSD9+SimF8+BIJoEnirkh+IJMtHn
tBpMhSAc+GBEnVbkVG2slS71a5jrThMFaXBwN5kZSgKRLrPophOBIpanTMxP7EzX
ito2y+cICH5E01aarulUK6OpNKsDEX1hl7QUCUEiMUOA5L/SGdt+XrJeFYxP8cn1
pZ2sdu3jTyXnElumXsCuJZf3PiFuDEEy/QwagnPIkR4d6pFMi+tmIztoomJIXZCk
exQYTZuiLZ1834CDl2K241B82c9IXDLguCzT1YFl9IqZhnsWmMBs3qJVxkCZCBNM
meRt+7w+hO8nb9xHS5qNMvi0Yiey2TXknuxgo7IVaCLRDPdpUmpeft1xOvJBrVsr
R2dCUieVoUhc0uSAyMjsctI1PlOG3WrGZa+o09aFekWQA6uyREOqhNDs7tRXH1j+
3n7CnoeDq6BqR0DeWU53dmD3d1dtaktTtchhz27tDkAO8tKiAgAYeNJosFVmW3Fz
hbL656TT4BVhIKB9hmMFnLXYM9869AghYrFABBszgq9gZDMUBRlOiCglBjJZ38h3
GYQZEdC0VIKPlzLYUs7beYraUtdIDjldtnKTnjdm0FVNEX9a3b51KerY9OvCIfze
KlzJwLX6vzp4FiYGwfw8OhMxUsBhkYsFyt+uOQESSPMPjbvFHHGCOxtL/5244aFX
s6pkTX0egqisNnAcweDILH3uxzLgp2b8hZGGF38K1+Gi4miI3T3hvM+3a/Z063O0
KU9n8oJvCudsUJAb57ky8Cqd2+G8/S1jfV6r7wSjZizBJdcqNBev92aQcTV9/zZd
4fKuezXkry8I9DIxuodoV8M/YJYaW9tfEPQmzXkGbH7cr7AZhW5x6mFq0r5E3ms1
E3ZQpnaLqD/B8zQCL3eAlNcbI3BzHSGucFmZ+sEKGhc6+22iO0yWxWh3cGxEfOGh
ge+riKr53zGX5LhOAN4fhEzTAhO8eu1vtc8lYzgocfasuLLA89cTHinfpIOMpt6i
D+EVTwhOQSmFmKj8yw558/RBKrymdIRz15Ukvzt9KNamT27C974F02Oi7eiUWpvr
b0+V7F103cbbovRqAuiWgnKWEfVi6gFx0iqmUiL3rYWtMjKZpOo+VsxjLe9kcJ0w
7/Ccr9FzocQXqb6I/DtzOGo6r6nmu1/0rD8SbrA4/O/yy+vimUl2DROKETKktfIb
fXfRinUi7bHiEckneBkq4euTN4Y/j7utf2NJC4aOwhyUeUUWc4VYkCjvP/ESxey3
8MEvDQ8Z14ncuTawzOs7p//9sN8TiLEZjFetzxMA/T5WLxaPn5rK3CQuW2AqXaiQ
ELQ/7HmQimtQcvMHs6Zs6t+qOnNrPHoS3GaO7ZmJfj/NCeKKdTLdzgLJgrhEOoyj
IVaV/EJoznrm/cKefyH+jwsf3oEZPbxljL/DZAD2VhePwDCKd/4fPNwH0YyhuKyL
RwnvCmPrF1M8n/JkY3gijKYvYGm4/GOv2TL+Lv+66BxHCLf8Iw3qaXpqNUFEFHjY
Q+49s1Ndce/775CycTlqVCMRW1u66vZmnXgHdknEO2WYBRuS0xkrlcKNCn/BFGCx
m3uosu1jEUUwcjGux6jaVfMIM/fbGngWswnHwC1QKID8oxT+c5p9M1WQhTpiqsWJ
ZlTtLhirm+xypm0qbWPSoXghac90I7X8tg6jtLIclUGh+nVjzm8WK53hTNbsy2ed
eHyplB6ZxRzhXMnay0Pp2ToJxUbn3PD8+8vFohzoma2X3gJ/Hn0xGib3nGK0HqGA
NC9kegbpcE1RQJ73tSV9byD5a4rGRvXzRe8JQpIVhB4fw0Mje/R6tWTGJOVCMoT4
4Cex+0wKnSs8YdpBxYl7RiLsCFeWD5gAjvJmijk07fljZ2P+YDBoaMyXb3lWmg74
rpsyrmOrc1h/3iDrXfbh993jGU6pXqSXMgQC/l7S2Pb6j3VcuCxvCshpmRden9wN
lqYUNJHG0Gvqvk1tdw5qcSSmgxSq6ShmlpzjBGXniIKfjoe9kF6gzCSWICJe0KLV
8wOOT2MAth8Or0s4QG14m+fZ4rwX+dk+GRDjB5xi8Jj7E6TeN/qCDaYs9LbvplIj
pbtsXgzJgylzykiszva/FenYFG7Ju9J5Ere04/cGvO19dAMxNt0W/LlTId2/hHwG
1oA5f6JLymB27ZKK5tHpVibOL9qJHxCd9BjagLTIxf1MwRIKxXDPUuDYK+Z1t6Iv
aNxRUDfMIAhSw3c5NebK4yl0vg/xLeDOWFEJkWLNdO4M+XfgC8BjqVrULtFl9ed6
fkj3M0gE6mGPAy+6mq8IqxwfSRVHY1KGvrMz9dOz/waL75t/LZjZhW3qhoCp7aZY
W/t6JQdbXwpck8iQX4WImCYQN5PTluRqi9gg/p73ekGhIwdsBvcN/Tu3DOSKwoDz
3hXLt6G2bm2cQL1XEloNkJwSv2HlqhThrS3J6Z2dsv+i6zYyhsl2sVtIDrSlk6n0
ijb6RcHHDa8NIEmboVIrB2bLyoKsdEnIw+SETDZ2wyTcd2eatutJCSOzcOsHiosm
eFhZ2rOM9z91mMjY3MNAqeH6X9cX7n315a9F7c08QtRVgktiDwXXppOrRAe3BR1+
utsQfCChbCIhUbfoZYj8z453cgDZFF0KojEeq8rqrvkdAefbUZSxan9bA35LRxVB
wS56zK/BWnkj/v3EfgNNFyqBzp+yWRgQoXKvImXyGvlzJgNyPQ8Ba9VibHxJmpCY
dKdEeKm3K8oatMrJugVPdMxkzNbra9COV9Ivfp7joUvaGyu96LkCZBZAMJ8XoMJ4
MI+csvgcgMjzxqbeEfqqXZBiq5dimrryFKO3fTY+bUJNQpASf8eINJXed2xVIHtG
pjsggbtUgNnbwmm/xfCULPiW3Mk3edYjuPmCbGXvutDDmgxX4tyxmxUC9l2e4E53
35SR12+bkpA3iZqKtfExfmPS3Fmnl3VX5Qp4Lygg8L2yOudbfz2JxCB2OrXgF6vQ
pdQN95fE7Thg0rgjKrxQHc2OS4Fnw91XdBOyu9Ygr0gzQaLbBcczsfUuomL0wo4c
tSPUnqECs5Iqklm6leeTP4oKGaB3BiXh5oUWtGxRXQsLCSkuDkSRlZ4NtTRSY0Fv
zHSLwQy2+fHGnVz2sbX9tg2y7vw+J5xPJ7v/cb8M07iV6K9IbAXEwteIU23RLMJ/
upQUeVN7uRjko8fPPU79X2vjddRgcR1fhl5KzEgp/TZHb40eG5CFcHaooK/xsXfX
7dXtpCXzZhQqrmoeSX4oHM7+O+o/WPU7ESDVjsaTH734H5n7UMZcV6zBZfQ8lPXR
Rowmk2m5bWff9qvdf62+UuQpMtnLw36fIF6B9ZLwvhxhlTzInkshg/zBZToc4H1G
Vja8jiZ/gcBaWRE+1codCB4ycesksZIwL0QoiYdrSDGk4E/IVqbuga4YEKeADMst
vKpFqskTwlktex7LDwOcQs8miVMeB3ytifUmfPDlEjgDLX9Ktxfi5b2xlPvhPhsp
RSyiB86IFPaqNKWTZsrWe6T6DBEBbqV/hHBLZe4SRuPsrBNsVJefOQBpqsIHz4o/
qe99VXzARRiV+tFGHmXoH9u5h4rzoxfpQg1rltwNpJXlr1fOmZkh7jmAu4pdUpY3
TYhoitjKjw1yd6AUmS1pN6+EsPeSxPKIFHtIF88JUrkEPYPAihlicaeY7yNakDDR
4ggcDtSEpmRvf39b7aXqkRh38CrswYxREc/uy6R5zLjFboM76U2UA/IrvtIxWUS5
4W73FpSBIMxIPBmgZ3bT+y4OhgmcVzyk2e1YcNExeNu2A9WPBc4jn+3Ci9TXyyCU
gf7xHE+TJ9SCoMzaxHg8kKciJpLBmascZiMDkan1WA9xQs3V2rjySqb6JduqIuR3
w4cmrMOfj38G4lfzynLTg1j1dkdOSyeRGTPUvRse+Bct3U143f4bsp156MEu/mSM
yDXos3SH2Sf6Danl3yvmEc6St2/WEyiZ+o2AVL0YasvOcZWp1RScQufhMtIMDwBN
dqeznrUBY7hY7JkntilFvydfkOG31g6mvZGYzJq+1l1FWylq2Yuq0oZ1LO2RWGAq
2YGExRhZMnYrpayE3S2Ys6NWptrwicZxnA9HuTntrmS+XcGrrVbJ5mMfPATicg1W
UaotOaB7ViIMg7MTTISvln38651kUDO6bwgEUYRlqZCGZ4QTgJkdQJd7lHq85Jdq
Z0TOpGL88XqUwO5N1uej217FHhVmh0va3KIJfA62SRSJgDUBRjOirpM0DYoIsw+v
+T3XDTDuQq0P/JmcPG/PLfvbborEgxzlcc/7M5hQNcEckDSoM4amMwque6WX1JEA
GgAFcS6TxSK0ZUObUltFooFpNyne3BRvyR1Yjwwfp8g4DHxB8DH4m9XJZriV7n94
TG0HLiLyDVgEbpuFq95QcRXL/V+w0Fqy0Dhk3VhBDfXrWuQVm9Iv0O+CRmDJX0KO
LJQJxrire2wl+UdL7d32WmDl5GsM1SzY9BuLDg2EQDapM84t6mcXGa6j3qZJ9oRu
UMpHiQr7Jj1PNnGuReRGXSxH2jI1D8oU5vLOtBKe6BtvEqqp5oy0iJd/w+2mVUOF
8QsXep338ObgQJXNHIJe41rEyYzKUOuYLGcEmAvv2hx958oA0imVPp9YyxrKOgPw
LjSu248C9hhPYhC+Ytmb3nrFail4Pag8GT+3B0cuzsFML7lyKVeYGva+KW3iW0PS
X3rX4CGlLr0KrxrwxTZC2Vx1/Ze2BKK6eZq7YEmH5ciFF7DcmOTz4lCm9L87GdKB
zKuf5VWi9kIsZvv0/SFwndYLwPCuz+uLzVJujYuJjztrtivoX5uDP9kytw3u+tEO
uVmU29/PMZGycS28cIERSzFNeZ1j2wRNaqlSPmb2skhnW1AT6SRJTxXsFpvGonvg
Rv5P1MNEDV/QqoiFjYf3kD32mAkUQjRsv7NrNa+UFxgUmO1FBDH8fwAUx8u5DzJh
jBEw5WaPDhMRj6piec/DLrzNMYOgV/ciQ/AKYEgnO3aymhaa9/SuGRJ2XHV1+yvL
q+QF9Bi0RwkRox3B585nD+Dihf9VklDNMTP6JWD5yrEJDBN8RFygDvjahQsh08XQ
ki1XrKjUPKRYCkTa0z65MIroauVHWHRx1RtmodxEm2DlwWcalq+/Jlg7AMmciFs1
Hnyir8b9iveh5TBzpNZkBI6EOSa3Ql1MjGpritqYhWUsdO8y2+q5IoFLk3ddTRIN
t/hy9EdXxsEiVyRSeLAgTzD0eo54Htj4qaQk5dldHPXJ2NhsgY7pTdvpZGk/qCgK
BMDaOpalZIRZSPdi656mqk6zHSiyUUH2qCDYswURDRWkl9zmnP/MT83Bc9QsoPrb
37difmPDVXQWTdpMaTz2F8WRUr6GYdfGssAMqwtPOCGfBhoI6tEeCBVwR6FULsZp
SSkxBBi/w8FAwSpNP4Ec8s7m2a+mY1K1Y0dn0+npJXIkV6QnjFbyMJ9j1GckKsws
7jhzwHtGQKOL0eQFfWQVOa1pixQPmbOk0U0mjQK1mR2OgTIdqjWvc2eVf+WvMFmy
phKawfJW7J+L0dKvPAax2YldgJJvqQwUBoz4hhFi3diE0ndhAlwBSoHJfpoKE9N4
dvo4UPVap7xaImhgbYR0eWRgVPMNvyDNewBSZ/2zJDQ0iaHN8W7vZ9YYz5INDHBg
DOUAu6cxRq1dyDLCQyJDd6u1ReeYdem5N8oQw9VMCuJlRzRgyKje9mf1BjWXlbjZ
ME2eY4+e2Vx6EJnXiXSCr0TozWIGy2M50YS/49lRsAPB2Nt8Zj+4u85HfIlsmi1G
OoWdLv+qs7kzMrh0nwGtrW8s6VuyGFiUXqoPOBYqeyZg23xbSKD3dCguDVH90ZaI
oI86o+kJ/SNTM65YJOb2gPQ4eybH7s7YWGAdZwEtbQOaKvltupc7kOaCiKKOzSu2
nXdqKLjiPyTxvRcGhl6faBjI49BNxYtlBTiOaNEmgt8ZOFjUXOJp8m3cx1ohbnMM
A68A3QrtvI32rfM8OnFGwGc2Hk/iMqfCykz5ZSo34ECxiNq6GTo1LL4mJT1TEkev
hwUxOZ0zGomP9e29/GQ13fTbCg5vUQDPXiTlisOKiPau5/9ggr/QLfmGiCU1tjM9
DVhYHRZRcrHFwu+TUqQHXRhVwhiHoIP6nt/LeEUJOIEhJc3wnSGJpZYe0r9PrKjy
BesKhR23IXz0W6z5jh2qYXmqGhyM4QNU/OwiGCkJWl+7LBKqNJ/DU3Bn2UjN+yJg
5+tskYocArh1h2FLPOLiXpr6/3zqVzveQruj9U4cwVfHlbF9qBx4XOpqhJ/DtT0p
tw1ah5FrGo8UllkBTJGwd7vfjCcU0ZnzYS00N3CuwmSG/NLQ1Q3CnOhU8Atjc628
HQTz9+AXUtOHrVLHkRGKi6SNN+YyKVFzwZZla+JTVq25tuaISrKbcvGDZAsYoH0N
Mp5FHAa79nmDse7lWhYnFUALrxwO6SwSg3jUCb4CQ8txUza8A/EcZA69lVnL/N75
mfBUeBG6yWTmao/R6vjAMvNRJ3qJk0mIijPGxCVtjlUMoe7eyoeECPUpMI9qhmki
wNFRfnjVwVygMiM5/crOeDOXbTM+ap8e4PSeMji266K71v2csloBVL2BUyALzpxn
Qtcu2YKBTgCbpM6BGb4fTnc48vgIM+o04mFF6BqAp/8dcR2Xq34y6qE2/MIBj7P5
pP6iTJI6I+bDya6fS5J2bN8ROulYlZn5HOCTdw5/QhGs7gjsx6bgHwtqVSYcnM5/
wj8mUrsm/S+OboGWxsPjKqvObtpkLSA5s/N4bbPaSY2l0D8oOjHtLWhtFGVEhHXH
1UwfHaReHFyXKTiWMTBs1iq7dqD+7yCkp/OW3zQdBRsycyDld7m9zIghJFTpIFRf
E9EMYIiu7HE7J2LR9NRg2/Gz4pws2cbp8A9RWTpI/YzPXfCxXQSE1b/1APre40rf
mkynAD63QzKbfmamf/bslxxJN8a42sdcKLfaVNUJqiglNInbmVMxrTRST2BLkMOF
XKhD1SeKGGvRUPDVuJ0pwHc5RdyEmmgkiL8JLI24SsPkcDQcM4MxiL8Dz+gqf6Us
9ZOLw73S823nd01IueAvjsOAFG4bev0NTnLsc/lIxGo5H28+LxMd4O/kzpvxCOQA
GNyIHO/SjHpoP/MEOhRus93AGeJ3X/WbaKSpeMvAeLR856Kr/792xz5jc8KSepxF
CNMZ5I/9Yi2GhCle5l01Q7fDCdcoAIL8pU5E2ReHoiMvtvkR+A2yWvj1A+P3uTI0
xCeaiNARJnuyg4IXZQzJjbr1hkcTQOGt5w2vD2kCndoJjluTN5N7KqlU1LRqYWnl
PEET+CYJlgxK5ZvuLOCUAKbgOWnXxKVtuP7Nmv7WQIInCI/i8dkk/G6a7DDTxa08
WlY/z3pMofIFNLfjd+5kVbP5vYKFPSQ9MP+57QoRWnrjBCcll17JYFY2zOdgNXXG
Prvwm0xrry0M65hB6z6YYmc0HxgJFo2MuVkRp9kfZ0qaYBgytNOdeqBMWzYnB2u/
LNy0Eiz/ED0zRwv2KV/NYmADGGo62lwzeyJurFWA0x/Dt1tmSjeSzFL+AkfckGTZ
Rn9f9TLoZlVbal+f2Bo6MYDfvOLbL19u3Z9LB82XWB82HFB+CWaRnmkku3bkOG6c
6polW3ggvO57U0Q3NjXViIm2l512CrSuxpoK80QDD6+WBhHVEfOUSXuhp8NBD19d
o45Vk1TsPenGgqB8xMnSmMmfOyRWoJH3rEkjG1U8bZ0Bjq+crNIw727TIyXWxl+W
Y/5/lZcQIBUE/bw1PVA4V0JP+IAM5SoKzLbcVQCbh7E7qW4S3dXKnwvcN7zR5oUf
6mboBSjxyFmlTSABGu+NqEySqGhzrTlz/UJqEdYEBUEZm0UWFX3WtZ8rou6EpkR1
4vdI53RV1IHhpckEHRJApZnPJI5dQqsKOBBLa8qwUZXxyt4lDrKGvCVjhoceEcDb
FKOUk/stlARRsT7ETO4OMSBqUvnJAGnNfUV7zska9iZN5488jdcZ6DlLBOuVMUE1
UVS4DheXA9JbUx/ebQooKVEKNhdFzPmPmiylXfOetnH/sJ8GCjnZ/4XWWg3QbR11
FijOeQfFoxlYPjEBT+ByYPgVPx/mbP/j5PDb/n4/sU+pnMDHbpr5ftV/5Tm0Ie15
fygQRn2pozhyXKB4gsqlk5OX8zOSjW5LUhnge4uNI6V0BNvKzs3ASfenHNXCzw2E
Am3MRM+NqUx/UAQlXQlYGWUwQ570XJTxSON1vWR1ZXVNtc2ZXJmMGNORnXw0ElKm
4cjqBemXGO7hWL1v0zkMEK7x9CiqJOOC5DJ2gBwbpNa4b+zrMUKbs5GzkKdlPFag
5gshiX9Tgff97CoSAMDE2dOwaznpfr5GN5j/D2YTb2ySyc6U/ZbCGEvC3tPhluIG
1Ee9099tCF+OvG0WPNiBoMfyiwazz1GfRl/qSHMe2HRuFR1WZCIhZaETt/uBrz3M
t13pGcTa5pYyluvE17q4NgFI72tBGu8gvJRRzfDVIXh9dsK32zWgCkVKBfBDGNDN
/InGm0QVPIY3WyD40vWAXIxDiUPtTdrqgf0qLvxEr2lsShIqKe2W4Lpuo++uh7xx
ogpGhIAqB1XD4p/lUPMoobDsMHxf9qoJXS0h8FqGr0V4Y4HvYmRBAXFMohI7SN+u
FCRRM8OuUmR4S9BPGWNTlVPoTf6IwPmrr1Cnbn2NDXOLOmHFCuuL29dAcstdtGZU
BclG8bm2OGUGQpyTEmSkFo7UwRzDv5h8jfsCPGJz+JNELeT7/vGZ8oR1IZMVOlrG
f/Z83AY2bSQThucmLmyaBoGinRppkULgvI2DD6vlK4InZ1Zj7T5UJtrHtb+R34px
3fd4DJGC6pP1D2VomX3YcbUYYYOvuIy/8VKRKsljGhNDFziY32jZezw2pl31sfa2
ZvXlufwNEqS7i9OPj8d+GOhWAoebYaXRqlqgHuFIqhmvchrnWwWc9pNB/19nBvND
BZVFAriP9OThz4Spyjkfng7/mH78IbFy/OHqdXVDMiC1bCBn2qgfiSX6/4KJT3yf
+KkitJdfZMrmhBpEebpHZ5BZT5xYYe8aD0zMLuWeYlyXrybVg6r5fjWhWCt4hr4c
/LjdcfTgc+0vusNzcuumq2ciDhvyMfpN+dXs0H5GrYT9qdnpy3IrQE8vE1n13Sbv
Wz7ZoW1ge7GZh3oiNXD9EBdtZD9vng0QlWlEcrkWZzX6vmOtK448jORGxDXzPaPe
mdnvBK5XzEcST3Oh+oOFqDjL0o8ST9KXQwcte6D4qJSCB/QHk8Vaohx+ZW8Wo87d
FQ+ouNz26Tg2IKhgqVkGizrtbUH2AGAi+65dHPTU+BXRpIl7pG+oxpy7uketQkfo
5XCoMOxsQJRYtCk1e20OPiPe+UKr5P2yvS3yjBvG/k/0cXIS8/j/+pI4eH0VWEep
c2xd88pN/xZeeq47n7W+Zq6I/idolL3azfE2C8jwKyyb5p88Lnp8oRU5ls+NjLpD
PhZEMjuBGWNMuM+dQIKd8X2UY59451S4h1YFnF9vwL91DUmio80EAoxyPiJDlF2h
dkbx2b83GClxIVR5CnB845oi4r2nKdXzghxmiiGYtTF/SYXc3/cPt0fvpPDK9N3Y
wt2UhyX/gPhzEZPOW1tXmXnmmcnOfaS6Me0w5cKtCqno/dzdYcyABCGNCs2vyeM/
S2G7sZ8IVQfhkWzkRYny5MecKYc+pIWKsmiOAlkCIsqI2m+mIy5Q5MeRp0J7Z9Gh
T+8DbTRH34Z1ER3b7mLKUnOxlX/u3VDD0Hxmolvw+bf5pSB/MEELtD9v3nfXEqpE
PqZpLv/lzjPUppQZdVFrX2qy56rW7hu2JrY8Bw4cbid2qJ/FdAxip/wfLjbKNn37
o5zDp9tgDNlk+VbZLCgNn3ApO+mghQ+hBX6agNm5dyymQS2EuRtTXswF1hkuP/VN
mqLw0VkROtJFHkjCZifdAH79lWy5WYuPblVF6hQC+74PN/xJnKvQZJBVXmwDRZMr
ORrNl4IdTkSBLiEs2mDqvG2dI5AdrjQ7fvP7HYm5WLKmy/NyOLIKPnRBMY+tv13c
C98GzBMhZYt2DMfQNTa3fMocCgkHuITzSH0RpRbywb9bmCcc1dtbiQrnJh155Yo4
cHlUKYRdMHq8E5xZCE5n5dVbhFcNPko9ShY41Kc8QM/HONRsFuDcR+D4sTuQ+iCW
XhrL2kmxv0F8f16vyeDDC5u6eHtm7NNxElt9mWj3agzzYB1O7nCGi/Vh7+wWpAT/
5bgw1CRJiOm5KgTP+t7WYSQopNX6UF7ZywwKLPXPgXb3GDNVCAHSh1/7fMizvSq+
LyEsDCbgQBht1zFdYaNt8llk65aa3wRcBVMeDKybLKQp95c4xpiTexSGenbIudsB
Aag9S46Ox1KiZnqe1app/Hi3nCAr5BbgRuttnCLjYEXmFT/AmdVGUdmVLSfhj/Q/
9NqbDbehqeGF+pOgbfbBY6tjlmAgahanYfS58lHdUXMSXMhiIDO9coabwEGZySxA
i+dWxt5M6ot+8fy8jclDc7TkyQ3YpyXuRI/I3ZXza0gSIM2QdpyPErBEAmZNPa3V
cm0tw/VyZyZVR0VvGPGNChVBliX7wvgH6SxvLOoAtKPPeSSeC/b1Qq99cTelcM5S
unMwYrDfsj4cssxE8D0ZGc/vf4mjxV0LLJC43p6zFGh5b/i9gda15YA8PPvX8tEp
pw5/iy2F5MIJ49J3w2QXO59820paiMrN1Fa59CAV3tEWXZIgT4vgEwNmWw0h4qly
16RJC0V/eaZeAMJbyLURMzlduYkc4GxrstN6XOBjO8AdDeCO0Ht9dhdtYlWndOHI
D+VfF3Bq+8hvLmRbVLsm225UR5kXIuH8Z/nHK05qJh9uj0x8xfwTS0dPclb1M/9j
Rf2/lgJuAqF4n0vzx/gAdgHPF5dVH/F9JIaheK2tYEZWZL5eZMdLfSmuxbk305Zq
IwN4lUiJhleti8bg+vcGYI4KHMPe26FAEDiuCI06lMiM/diWWkXXoGH4uoiCxe5W
lvo0CqmAdmJXG6wk+h6FQGBwadii0buFFF4/kERJrnpJ1FxTQxiZPQHYzikmi8Gd
FGO/TLg+dD85B4P2cqkyIkXQVMaU7iyYy3DGCg64FVlqSAu+WKnY7lkc3Y8STKl6
TDyr3UdZeGy5EVXnFNQfqPXoBatS0OetI3mivN2r54xShlPI1TaCzWIRY3t2GMm6
L1SKVVrUkgErd2JXZQb+DrhLhZgnabZ0NVQoLT+ZljOsiJWtRteKVBQnKClKPOY3
1GVj88SVboZIPslLXt1YjwhGpE4mf1tIGlrJfPeqwYUAUHwdDt1D7qaz0yFWu/5w
W2GtmzJVfDbOXbNU2EpICUoJuJ4kTCDC4phui5B3/GTvFHBV8tcwH3M7lbo45NYH
8+oNBXaxzze0TTu6PqQauti9NdVNGwXL1qvJWphX4R55Gw3J769OCewhZvbfvkGl
ORmA+mzcujgyLF8hPUvVY87RQbqNg3taLS0BMlyWj6yJmy6w3QeISMjBlrcYnvGI
vVhSqlPtawT9II5BC8njdLLqXJrOIfphPnZYz5J/Vl8okehr0Xa4zqCer46KIb7Y
8vM4kZK0Pia1vmkT0pFBwpjsvpaMIQYs2w4h6HlasWpo4SPUFMJ/Gilo9u5dcfs3
+KGk50sJlMt0sUx9IUJEeo2qSFJ32Uqm5yg3ltZlGywDaueYAmvh2C+dqiUNe0zW
CwhjdvJQ4G1vu+GTbAdsCVpk9E3wYLBLbQXwUeaQkuWPqX7rtDIqoHCPl4k/GHyf
aKJMbvxwMgAMC+KUD69yGOoKQ+D/Ehu9D6FUUd8Miwwu55rUpkpP3PLHj/uSJIOx
3f/LjumTTbf3nQGj5CQvfGGicfGL1RCXX4lKdJIpNWDCBEYFqlYHLSXq/ZZThEmp
bWhvmz9fq+WiU6qXXZaimid67icYcUhjF3+3Fs3TzI5czluyunWcIkAf961b3XFY
ldSTkVurWFpsepH7tB9PGs4wFwYifpxzqEmAdNZixIA7ezWkPfPn91q+8dboFMV2
me9kDWwPrykj1mWaSSSSz5A2aj2J8HDSHiaSBlg7ktmO5I2JnmAmmIOAYa17r8eH
77Z7r2piuzynpVTr31DKUNUpVLUFisao5ttIudlbA9bJV/68A0eA+lgbgEEV/U2R
ffPED5oOFLupYXRvqebgj4iRed8n4A2q/dERNP9+cv3vQrpVK6pR1tqpA9JCMlMi
ezJ/j+u4cu5qVpBHnJ8IINtuYnZdbMR3m7FQ5icbXef8W5Y8sV3RCmzKKhoCSYpc
MYiCrYupkhkdZD5xg0hIa6cqGoyFCGixf2SqetaXSsrwxKLZpd2PuHp2jExEaf+U
cjd7B1powBTSdj2GvM0kF62JH+SUQuzhJwidq8eykkuCiFV5pSd/DD6djLzfTFYY
+8H124PCwq1qh5jX649poSwGhXihpfVSMhirwSAwh2twNyhlEPjla54zp27kZlUx
23NurSRk/HBe5MB6nPyHjsOvbNitVQYWD/h8GSMlcqFfvFe6JvJvABeMZjsRW2S6
JLPtfN4RM1PDnfeMHGDVtY2NiHBd5w1FM3kOb5CuqMDzTtgNPMQdTnQe7nE5qWBi
KfINB/sH+vUYJUqrYmqjGIFIKdRnHInOum1a3E6Fu1+4CrpHH+0Hjk0/SKDL1zG9
6vuUEEe1w1LepsBpmkHfuKeyjJirNOjmgkHd2MYHTDSmO4XS76eouYVGh4GsJYoS
ZY2CHi10BLHULt4BHi9yLTAMlIoQxTRKPMtddvWhe3DBftY3YMxldJf04+/j2s0z
kijSNMJh4Gpag/BtRZgbAiHdZxhAbxPyJQ4WeLm1keEcG8LHPSYYrzA2YdUoRS9u
CYifZGZjja98c6RFYOYhIyyQpz1okPsazT6U5IdV1ZyGJ09OTlwh6Aw53RGJ/Cel
Qb1npbgH30c3wct38MbzwO40UpR5IqRUpxGbnXpweHdSL+uzrbiPEAi8f20T0Z0s
wDFSB6wdg7O4afxVx/XoSALPow+wGD0xu+Kl5oFafqmF8XhVw+SEPxXTrltbO55M
1RsB1LEYTNzXSAWyuJ+sgMiIA3AMLkERx6zSWQes3yNZ0pyDFYy4AnrP/Ru0VeLY
t2npH0ed1LeXPprMq3B9W/Kv6CBmCcpvmS57LGZvOynIQv2YwFtAmwCkdtTpWMvx
AeAW13Syxf4ORb6ZKX84Ap5m+FQ+vBXakqOCz22QD5BIsIt7KNmQMra8dimoWQhY
wcOf7R5Q7uOSSecGmdplZiRbDzbcdNYMa1sTM0hE6SlMzRdFcQchPnYmCmVmonbb
CyIVTCUXf9OxUtvy3gU7nIdRdkHCayHUl3m3Exnd+ryX6RH+BIs9KowwVzig/oq0
jQA2sai7NQdOT9ZzITJz10BXDotSbUEMwEQPn30Ibk+QUYKGA5p54ZmsnbmTrG5t
dwYBZQl/vqgnLo9nBiTqpwWKlXcuaYcowVxkOSt6qYMyibkpsULAD16jxEb36myG
FvrKK8N7lVIYNe3fKTCDow6dL5FPegRacqGxdRhZ1T0MJzICbhWeDqQopmaTLtmk
16Tx5ESQGxJTFJ4bFw1d3GMcXVbV6RhYNXnf2T1V+vz0fXMoBGwa5slK58SVQ6ol
aMnP9HZW8PuyIFh+ABU+ukKt1CzWEnytpLxB9Bu6cUPLawoJXzoZmzlpntPUxSi/
7ZltGz3ddh6/1pbMMBB8oo96pDWpwfQwKJ0emgSBlkB7IU/LA9ktCbdfBk0Gkp7P
OcEpBfiwn4JshfX6V3NxLuEhhX2fpz7SQZn4sMT/b9QP6Cm7ogXUB2zfA+jk53E4
gSo7zGVWODzO4+65RfA4kPb6bs4vYy3ECkuEc3Owpey+v0FBJMETcaHSi71IbXDf
30vfOQjbWdNWkydv+KsAcPMj28eR4GHbyU12miaNpqocgPagC3s0twGkfH4Fa9bU
+f0eltyOSAVuuZzJwJcsD8NokUULZHZShcRFOH+HV4XzytKLtEomACIQhx33P052
IhKj3+8TXoT7b0Vcq0Qiz+y22H8adnw53Fp9uecsnczK00rm6sEXSRvraNKs87Wo
/JbcxTBnz6fkL+F7CSZKcV/GO06+D9zOmgwS82c4t8Pf/PpvR5h9LOXgpKzgBjyL
keJuPuU1+X37mSqB/jiOPUNxXZFCVoxNCWIgHksWsypPPgpL/KN+JJMMRVvyXAV6
5U7B2CbOLgHOFQEqZwLYZHHYQW+u4hpRkYCyMKR8/IZ+JnkrhizyM5s8XBhGgF2t
+dU2FJxo5c1QT+Uv7/gjRI43ZCdbhUwYER6K3hjp8/s5xfKrHhqaZ1797TyqTC56
JOHuwHW0vZzkwmR1gW4uga+X3i191fo1LeS/2OPDf9ixvovUDV2e+MOf9W7SQFN1
gQ1+KkLRLNyxoyNhqeWJxPahTQCa3/yC/re6+mV9U5uz/mLY2aWFxmcL6IHckuRF
6hqyqjM8FJMs53k1wIU5gJqoOKMdwlxuAJ3qRkgyY1oBDhQ4ENIASWjNMGdRau5c
VQo/XcytlQTmtTx4rLLSBKb2hRXQ0eR7eVDnIT7wXuCNDgVhFKyf9d0smNBd7gbj
YoyJ9aC9rmIFp4NEogTblGoPDMG/deibx+nJeGWzgt+Vwm+k4vcmEloxXdQGnVaz
CUIQzwPvMV0MYdUC6UFDeWyyrqB5m9sDQq6bcBYrwxVUJbLCKr4cAoQHzr11mYaS
HneM/eonbkvpqlcmdALIQuMGJaSKpUnnA3SZmQ7Ib6JJaE5ssk5H8ccHuifVlSGK
4xDtz4I4Es7t1xzY8bp6swPfDqGJl3Dl0Blbk9cSokUXf+rz+64XgvVjsw8h01zx
EdODUVeKlh5V19VsZ1H7GJVc7wZdTGRhKtmM8izkO82hLqpuIEK42tcp0IMRxO3L
NAqrIgnavACUWv8zHSaQyKlsTLZza2ZBfy+XuwOSmwafjL9dmak0GwdA4ETecvcg
urq3Pf6StbcmUZKUfQgecPfdyb0fhAo7klRlk63G1HTFYPYgyoJt/rNf/n1s8Liq
T4HUJaOGEfrIcxs3XipJkSgIz3h0fMsMYO2IipedQbrE9O15schEiJ6SfXXpfE3D
IOL3kBg2eb5ETS6utI/r6KsWmk/Ov40zFimVb3wT0T5Mn5FY1Tg1wc3VTztoBsVC
0oWYEGy5fLMnso6YF2Ww+Xh9F/hYqYgvD/e0jCjvOea1e4BFtll4kTHdtLhI06Ve
cPvweBwckddvrmtXUnc7HkeXK7tk3de7GK9/ybD2olIOlMA0w3lLq5Ct+TEm3V2a
YamRI9ExywH4816wWgReNI3kFKVms0gy322iYgLaB8f6nzOdM+vZyembfsFdoCua
+KKqOVBE9V9fzwfBrPo3AWWIZSgFyAm83W819dK3faBsp8HmQSM4t/9vecGDAtfc
sg5S8sH+viXmjyjpR2uQpuOuzVbgX5Kl/N/Q9/x8CLsKfbsWmSsIRMgYGD6liliE
ppT0NgyY9vG7wrmv/VbaS9XXx3O/llgP/OeiwNnP8l9Q44G+RBK0nuqAk8P6DboM
G66wneP6NW6FSdAVWTbygQkiSO69zbBN/RtGjHfRLemNA08FyboJnQIzVoJUgbSS
gmY2ihK4ZqnWcpO8XiKjD9AWuKGL5R2NVUvwu3THDoS7124dJZuql6s+MYw0VeOR
d61Q70dhhnkQY0B27f0Oa5tctcDDDXRSxrmUY3dvqpO2jyi4c6sEiddRtHe2WNHN
atfY0dwLylJnJHHDNsyA+Fkhy8+cIln91WOcaxlVARgdY7e8q4u4w6UxDRDty6eo
z7lC8Q8ibJ19BZli4FwGi00afns1xtXNVQSnVR1me1TbmzHt4TdUN62R314mPrCU
7JjsUEB/wy55qUx1vYwsrs1M3iSm13NkE5VlSC9XxhO6U8ilbEGacUg3zGLQWCrV
bl+8gmhzPm9PbU/l8q8kwrqDWq2Mv2IiWHWcaHp+FTcY7mrojC8sJ+/dfyaR+cI0
+Zl34ra08/smvuB3X/IrQOiApYtke9B74ot0kCr/d1hj4Nu4W/24jc0D9+KD7d9z
uOPlWha7RE9zwY+rZv2kjg6ToyVHAJN8f9hb9Lc4FYsF5ooW0lCrf6/kvGdWFFjq
5+4KYO+/mB6tAkPlYsLeEgwFcQ020H5EXhLmygumDCRmfKrfl82TgY9wdyniOMcC
A9V3vPMHwet5jw+5dZiBlEaSZh+6KGytnyw/UQ68pts4a65k/PtfDbj7BM5zphxO
+sst2B4qoz/wmLXYzgklr47Hr/gHG80H78uYvXLnYjNt52s9tgvpYxj99/H/qqEL
5704sRAcfU4URhCaX1/5DSXGCML1zHtEZqQ6s2z+Wdc6ZMGoo6KEaRSh8yn1Smjd
H79s1NBoLlNnEAWPJATYIvcQ724xinL90DLTR/OOrFmf9BDqPZOpD043uNT5Ax29
s/yFb1ANirZWf1n219xkY/L29C/aBao6AM31metmTxXbgi4rQCEdz8SN/DecQYNS
eb5+Qz1Mv4TcUo3e1otJNMQKHG5rrKU/NuuMMgehgAgqjXMX53/LcvGBtFjw0HAM
SvfReWCgTC09FbOTzTs0anKJSXWiAIeaJlYMAQZCpMBwEL51rg6czRIBEcCTH/dK
/a2z6WqEc9KyoOuLd/FwK1HNmV7u3ELN0L3bEDaEdIZeDbZk+DpWl6BLPgp6ImVa
P81wre33rfVRn2O4XMUE4R61OXYW70O4xLQ0xoD92izG7DweyIUHCEO7+Rk/DKJf
ITlr1MYfmqGWQT6gOknIDQV5Ek51w3rerBu6uZqkSnDM4qMd24h73aEz6ffqdeRe
c2bJibfjRVCU5je9Y3OUDmQDC6Sx8AsHbr7TDo4yvo910KctxesUepCnYiPjtgWL
5mZuNldnUeugVQVNf3+1unTon1tvjQtPJYrCcMn49l+6tVkLd7gaQuGbALrr04NH
kLXSSe3Vt6eXpMFntC4oLparxwXZ3hF3lrgROZRafB9+nrThWOv3h6zMy0kn7eOd
n11rW9DggU5zSXOhsqLZq++A7k4h00ggKG3JtX2ukvqbsVaBIEdLIyYOySrgzVc4
7NGTOpkcTNsqC7wJ0LvhPZ0Mjn5c4Y9UeFRoC6XOdK9yFXhiPyTxM4R/fDUY/n5J
U1zzQYuvohTUEV85VtSvpeSZYmNZHEbMiMNDdePtBcN2tcRgJ6LgvCA8OugYUW3I
Azgy2b7rfqO/XIQe1BLYBcsPrCyyFUPT6JiDW/ng0yxkOmkwR2nD0qPC3K/g3AAV
3LdbC2Qv/TqxO8o9LlwyynvezOEjFsxjh+a8JIxgy4jiHKUhfku1k4iVW+ESAxRn
fi9X3yl8o7RD59ghnUJMOmjsyN8m9iGP+iChcKDK7OArGH5PdZNsQPUX7J7h2IOk
O1boDPW3EaN1XQ/2kQMj+puV2/esqQGsGB3645J1V3HfJxkua03EvEP9reGj/d0E
PKkyOHxdBr4LS2ems/UcjUJlolwotvGju5x1cZZq3eEqi7aeTAEHE56JI5KdyR/U
GsafiUhDLBGMOBIVLCfA9kTzUdHFcYXPlsnJjecazLhqJxTIbQswEjR+SO+krpU5
f8BQlw7V/J7kGBaS3IAfy1pAkMNeLTH9jRJCgBBdTjrdjjgeStaBq0139T6+tR37
25NdXc3WuPRTFdEfkjZCnemaYbPbE2o6BsRylQql+lBikckzZT310qRlksuoTdkC
EXyO3utQsbQ6WUVJ65SQOpSFrVnfExtd0jEetIyga31R0bn5DFcuDbXSD6fGJpcy
a/Zmweb4dQUYKUvIc7TX5JtLcqChKI9SKJ6lLOoimbphXQyETZBdo4CCJNbkKMPg
CmQpnqiUXJoI2LemfyuQB/kPc4dE3elNdUDDVfjlNGZ97Cjk9GU2I1SAuFKEdUOq
+ZPnKGE4w9N5Wj2pbv+448mfL4Vz74gFXe13w3XPNn8G2ES6drLkDDJtrYY3qxOO
sfJhRbxDzZi1QXbWaOitXzgbgCbXYYdbb7g6BKXKolWiquynm6/ubZv3gkgTWNvk
4dtuh5o9udpwo/nnOF1IS1yBQvAKxNjSQLtv7HBAHjNeFX81VwK9lkBGBsQCZoNG
Y54Kskxwckg89m7IvmgdgGHKk06FlRyCIeQnyxQHMjfK8evl3oY9IRIxC6Zqq8Zc
Tsz2cmsaz7PNWL/UmpXVL/0ce3NjqchwU1U4qaDGqYZoEa5ZtCAPW3mwGFyt6J2q
pHc5TntdSGqr6czrMfwuBr5E3LunDXSkknIkZhFTA9vkJF5f0/uFc1OB2Re0wB/O
ODyChDZPKVl19F0vYof60vbBYcvO3B7fEhGazuiaNXVCyC/a46l5xL8zxohzxbid
3KPjpNdArTlfeHWWEQiiT+HqSd23QmVGyEIFjcm5a0JqbDZk1ao+VQeDgvB+fsuV
qUcJmGcVE54hzq3JCEk3hUe1bfOFxaoTFRWuV6yKdNvl7hzoTnhEsr7ujNnQTruz
MIyZdXYAu0tHcVGqKKKPHwCYCjs+JBYYzBlGAmgLw6ur7FLs1dfPZ+fWfTQHRZGV
B5PZDVKH/dT642OwQDmhLKgy40DBJDZlh7ItgOKv2nThX3vVr7codsflGDwR474K
WD6TojDybRt2kxtaI7ZHRKchhLeyIzaQMboWoNLC8XyAOUxYlYM0weUGX6F58SSD
tu6JnGJwbvOw+ZL8FHmG/dODu78HoYmMT7eNX1OBnDqbqA/knxa2Ax6OCk+sCRyK
Hq1YWTYRnoOV50vtbAFXNF/39dxoG2a2JtS8U/KM7bkrYqhxSf5lKcTfipbIIueW
kByOh7oGX9yoj/6/bKzdmoIYmr23gOebm0rk00+aW4Brkwywg9hf/jnw5WMPCP7e
1i6VD5/Ldh/PChoQZ6pYOhSHps1TETuvqFZhI8kZF15WCOu4//+K5tSX8C39dB+L
lMNJZfBmGOkdgpC1i3VOJevgQTcizcguD1Mn1bE13u0mr8zYc9RZXMIQ545TOVff
yRx48SbjaIOo6ewuxNk7aA2hA/ZqLC+Yig/zBdvxr2B5zWiCqrcJ2ytV+cDPdvgy
fhVB7HiMqkU0ArR/4C8KIIbtIumWM0umQiVIjXn0qKOn0Du8VSt+IZmjxfEQnSq5
i1u0aeDHIHQI6aT+9jhAdTzGwlFJHQd/GVQV63CesAOnvULTvHx3yMTjINWNf79d
IPMEiDo5DWHDDesn4OHU7ZRUGRx+ij2SDaJBREWEt4VXqxEBtFpfEqQ6fgG+ImUW
PpquMiAwP3aO5QF+5v4MnlL01G2U2wo4xhxJzO/j+Ig+60M6SFrD1RlWL4B+I+wA
wkPf0qUBZP6WkS9SvR3DA0KiDWp3Ho6+OYxHXwzVo8RCTIcVsGtXH04/8vhrZDAo
p27bVov/w4OwjzHU3ISSj6FStN9SwBr6JHxZqTntHf5BcqVILNRJGyF3uni5qyXv
MVBl8wv7AJbSffy+fHLIxpWyetXiF0rOq2zY/7aq/cmX7kGKT18yHX5fAxoB+ykr
MU/UdM/Rq/w5iT/kyeGO4h+pvMk7ndaPXFMN8PfrMaSwC4ZbBTEQuvlsO2fxHRY1
XkJ7bk+/VbEI4VJ9AHpPjh9D+D/McNkPJ1uKez5sGO9uWbqI7gqGoxV/LomD8Rdq
LKROHdqOTF8FFUc6H8mYnNVQ8yk+LWYRUsA+7cC7Tf7MteRpN1uXoiv3LSy+eri3
3+hB4aKEd7ZAFa3tEYFC9zl8atShQ5eR4Aq+2PhB0YckMyWcVx92BJo7v+/YgRKR
IAoaDdtAGdBlHBK11q+t8zFLbZUmwhkYOEY7LZKihhITx3UX7RHkn2xK7282woE+
CzVom1+bhLhW4fjAHAX3JMm41I6Ys3CjVDoAAbcnheH1Fk2uznc3bgqOk+B5lIvp
o000qjAGs54Ydg/0UZB+Fj2BSq/jg7DNVkQUvW6HFaju5S3yvloBa3evhTCFJLuZ
qH767Ffq6Bce7IU3y20z+POL1k1Jf2bGqIZT3KxJYS8ug8r76JY6xfKWFHjXfyIj
gAS8aSFkpmx0KUJjm+Qyqs1wSpPJVNUUUP5pm2AWyEEH3O248Ap9Cu6Cxn3A7wCZ
mxYue1/88rz5iQYfzez7st21fhq14+w1VFQ0ZwQfcEqsuMu9RcOUqUIY5a0eChpQ
FZcQCfSTB9BfnUTM5mx1eV9pIHJaW5BGlCgMs7Tzz+yO6aIYsXUPINj9H6uRtjY+
3uUrE+bLkyjTRC0RH0uhwCkYIJYx9Pg/V9iECY/zazWNDBb9GJXZpJEnv/8Xx1Mz
5NluZXBrOQuMd2QlxvVuafutw+wTh9DPTLVJbjaiYKF59FM1SQteRwVbg06CB2+c
DK2csGbLsPea8QQP+XUmioTI+rkfiTJ2CDL1ky1XJykdZJ/i34yzM3yNsJSTgxVb
kfzvNQ3vHhxz8Zho9jD9MPXTbLn+CzswyuqYqXFSR0jESxCYv+gcKvspS0rxnjgW
7lVrdKNt+ivxozARRhmif4cJQu80Ps8vK1hOhjo3kT8Xvs1+Bd9XcsG0Sgas2jZk
dsNw4UgxYKaGwLF0+oRbCvggCVXjtrn5ViWqXQu1K4K1OzRfffnpHSUM/HiGsY4y
EyIEy584AW2PG98IXULzsuuqpw+jIDool5x2gu6NkUYybuRsTW+ZPOX78007pJ0q
5Erm63TPGp/yHqRaPVtB8DWVOgzCC8Svzj3NA67C3dL/asZGc06YohfZW11kbAlX
CVVzQXy3+96w7e6UKbZ20khrAgjwSFOgde89rkZGonB1rOZAzG1bBU54hqN4XDk+
VdiH7H5H5dzIWIt4N5oXyW7uDP4BFAgUIU09d1FIEd92Y4L7ur0ZPmMF9wgIj1UL
hrhEfP3EfOpaC1EGBGaNuc9P//ADY8p2h2/blFiRxlgEwaqyWcvrp/QEAnIJkgSk
Up7tsht59/w1Hj3qROkSvbSn7EH/5bAvbNFsGtK9Zevt2lLEEPum/WoD/b6ffRhA
al3umpvpbcK2R8kV2BMwbEzcGUV5elc+MvVlD1mTA5+/GODgtUeLbQGziksBYfnC
0m09LtrvDVceMQxQbmsw2WjxYgmb4vwiDosRrVSXVCjRYpCTgGiap72CPfdl5EgD
JgHxw5IEVp1Kha1kNItZSI/bAMo3zlDNnP9yUazugbGDESFClDE38N6ptE8gv1nr
AqWsnleAJT5QvudxAONIuVpEncPVjydjp/KdMBntQAejX7Q3ij/02FNDsZbAVNZw
zzgpg8rVN+ozR3+3wpuyqmjNCAD5YDyR1tSd3zB208xCJxHJowMA3YJeAj6PYar3
zh5rJOV6AD4sY2x7SzG8eYafd51rI83q2rcZLd0WmYn8gMeL53oTfXTRcCJO67Ax
mmMDb/KgMRvv9iR8jXm3iJyh+LqlECiHHJS5ur0v2YSVz4VzKwcpFUpCj4SqZSVq
0uUr2BLTwMWcy0ARw/uHa5ndEz+cqFqTi91PQdpCLj11pz4+Y2HF6mE5BqY3ooMH
fbj8/nrfD9OfWXfXfLZNjayVPW23VxsWJdulenmjK9wvCSoLm22JQ5Exf/ahGCKq
xuWVwrHzMoZZhFwdZ2/IN4HMy6PCBzvNiXDOzOvjNVjGzwhqKpLw39An9AQBaDvp
2LMc2Jm7ogYILUYGFtBZZSysWaI1HaSugdeV8qIhNJ8Si6MsbY5/ctl8HhuTNRuc
fUnNI4V1k5BNPJTuH4fkEgG1OqyXDfJ5GcWAJe/RMQOR1IHlJsi7xz+08xeXBpBl
ANGKzjzUpmQPp+Ld4uYiXV08DhVNyNn8z/SpzeCutVhU7n4AqZoqyeHHqyILGslt
pT9eod3fyTqm+e9W0Mdih/oN38dJrMaZ+kNXpB3aXgedZF+p0/sf2ndDuFEkWHaT
WQNNW5Iqu/rGovgZz0xl31qd1lim9n+Fmfng3GX28o3OB0CQch0gEIXmhGnZLFE7
jZlIHeDSrT1QL9QjS2hLvpJanOXBHMX8whwqWrJ3airHyk1B8jAxFtMgfjHlwrpu
QDWDM4geSi3X1wg6PFuqbhRhbxuDNy2snB7jv6AMrg3rC86Kua+B+PpWKg8oEA6t
rHxK6RA9bALhaPzKZtkCaB8vJGeXmH3ywOVr1/uiyNq5XFhWOPadSK+ANlO8BzcW
vExiyQsOlJbJkxnBwWXzxnvpDoSYCuc8zs8C1zJt0i+YmTuuqWsIwbtcyF6wr/Cc
JX9svZsRxGSx5HmjwoMLI+6xF+nGx1gFK4Dv3oJnwA/SEwB92LY2PKQ3UG3OM9K0
WlrFJJlw9nbRNdVzmt9e0tB5ugmIvzwuTxRzOWVTB00r9I8+1JeMs1C0G507Gw+7
yh6Qi+ttEOT73JWzP62T7xWL6YEfVfdeoLOgyak+9jRr4L8J5ClI9g81b7SPhgAa
y+ZhDiou6/ipL+RXO96+AYdoYp1vnt9bx+aeZ59Tp6afFn2f/LmNCVuj8S69Mpbr
s/iXhzSwqRp1Pozd4Nyj3wiaOy3vkPyT7VikeFG3bNe3UEifTpzKxcA2OIt8hVkx
Sk4bOcb+A5VzXLhdkBsH9l54tSJNKYorj/GXbIBhrhQ0OtxnYL94LPkLjmmFl8Ll
prA07UK14K8KobqZu9f4RlwljevTXbh3L1Ik7gvS8JKT3eGFPXqiAPDxJCm4hBJ5
HxF3BuxQGC83ozHvkDqTdrHcpCgUfyBu49B0GIiOJm8BM5cjWxPCL9iOm78ANDKH
5DHb3kem5Q7a7zp2A301MKaHt/DhbckFlxUhYd85S1lmH63rsjH36lLJetKMe6dl
KhmvnVmSqXDG5MqMiYH/u+/Uus6rYG2oHKLi3a2bfCdsGAf02/p2pgbg8dw/t8oZ
UGl0D/W/U7PylROTYJfsc60gu+KNwmk2Sg+Aw8P22YQxUVUvs8xfVzAdIIEEv4H8
doSv1aDDgWBFujkN14VU8jv4jVs4oy7SLgaTATfXuyrbv6+4sJfTEoQZ9Galg0ag
+Q/rSWO8B16eNp42ZY860xrzsaiIbdqZERo9Y8YgZsNDUYv/ei2T3GTKgnPxrQri
v6vZhktEhWfE8FIPunnInXwVCUIYSoGyqrEzEjMl4MO2Rrw8Gs4y0QWmBjmf4d/X
eOlvdS76tFlyiGaPDM/G1RGyI1c5CexQ7ahlTy0+eC0VubKXEB1Z/5HLFsjnzyn9
PhCm9Sc59Qz8hB6wrJUfU8d8azDMnr2UF47J6OHF44b/t5E3K0QAN7Vp8kq/crba
B1KqHjXNSseYveKthgAThoxSDAtVACqD7k8+3L/zqCCHlX1LXPwYDEUsqJVlOrCe
NFj7FNHQ4fZcv3dWoRBN7xvx22l6M501glgLJcRnlO16GnqnI1PScvucU0Du1Hfg
6iNggzVv2RTDEtFLArPuabBNLRIfIDvctFyKH4owwoHhQ19vY2LvVo87VSmKUmiZ
vNEkPAvOkSrxXIEs10X5vRpZs58sUz/KNSkxhR9hJWZ3I66tA33hsTqVdQOa99nR
uzhma4UafjRMUHEyoFAQ6lXoS7lP35qsO5Gk058n8U2/RLIOqV6CfqOerS5ZJs3l
yr8p+jHTHxWOgxp6Rbqsu4OCucPnNx/Xs/qorqc5BJ0vRv9mVnElU4DN0pS5oVNP
GgrcU0fkdtfyA1JxDbCp4FjOFZU3GjII4wPqN0uI/9ijlNPVAJ4XRn9Q5qcsQRaI
ndVmajVkziQdC1BiFZJZh9bzi1qiNgcS4IwKNWqX4LlUQthAPeROu+58B7npy5av
Q4p/L2v3EIc0snGdnKub1/FmUtC8Gn2iya/tUvX+S1UCyebiWYwvSXgG54/mknKk
xJGcrKb8JdkESbf0K8LvR32nEqwD63k0kCCqyR3hGr6Ql1mwcJbwRG188sMEqNp2
QZSeZ557G4m78GV7Dy/jrUbAKjyUhdfxTar1CXS8YfFOdqpPK8DXuKfcvHN2mYPQ
b/4SstQlfvpcFtgB22iCvyCciluQLCIFQ8QZPvK2aFPhofZ9NbCW45/Sj4H4y2yv
5MIGSv7ZcbyrCl4C31VVg3doUuN72itbC/SyjHXLoOeQMNogWtX6sf2pjw3/ROvH
2TrMRDu9VPHd30CbrfyU5NoLluQpoIwcvOClpmoMGFrGsc35lXAWNKbN4DAuQ3VP
5hvkzE/Jnt8gb6O33GFJZIg4qx1XOZtgi6RMQ5vcbTFcM9vy/tFFz6zdMM+CcBLq
F3cn+J2z94ec3tx1zFe+Wlwpp+E+blt2wo+Y5XnOg6kp3p2ZfbTjwGPBnnolYr22
VbjD0KyVGsdm0C+5tYzr+G/4u3Dajim3f15CBlipa+YEHnMgBOQ4z1JBWJkegvtP
6moXx1IcPfOzM26WiArnsyPNTwlTRqLm28TpqWzdvjcJX7KML0kWoYD3vEfgj5SZ
mJ5i78VIS4BXOkLVnEMvIKu7Q7ty8rG1clpbN8AjeXl7+7L//OU1M7OMq0u0aqLh
HuxfkugzcXlW8C+iu3mqk7BcrWfCfzr75juDAJqvX0otA8Lsz4oun7mb8YNSKcyy
sYGqYi5kOmguVoSubEcLxR3cN3vONdI5cPhmZH80PX/6sNNI+l0CKhKlLXQxcaHg
r8XkJZ/EaiGpIxkaBs1ReKhcmZkWGi98IlDHtQgrwxWYukcXyl47wv3DwV7J8VP1
YMU8FOa8dlnkqLecVWwTLy+6EvnQ/wqY8Z+eb+yWvMSiOT4RLjPpaXBosO+alZAY
wnv3iSFnyeAOANjXiW9X4aV9qYipIJR3LIvTkKcC//YtCJYtzoG8Z/9Lt+LHLKvA
I7Tchkk1He5U0LS6zWHmrptWWdRK65H3js/yeE518t7tEmrIJIdFP9ziWRDMq30a
DkCgdEAqGm1VzSX0kQ47jMjqYPL3Y8oJZiFgDGLQ9oxzV8FblR2PvIIIvsf9igi1
hfvlRfH6YNqeiVOrTrf+ugMjI66eHKRd5dYrEyQjvw6DD/FyuNGxX7sFnr05h0F4
iwrIMJNykeI2GEEP3f9pDdz8OvfC9YHwtCuVhdUqCYG840nBbfUiGDNCt5TlNBp6
0JwEy5CCEKmfV4HZ+c63TUk/IlO5qsZ6g4lu/5wRyd59+tYYRm86jk5kRcVKWCbO
L8J9p3wiZ1wCluM3QMUuq3TcCCQKWP64Sc0pKDcY5liIjwcOBQy+y6DFhi+SUQSW
/ORkbJ4V2co/V5XXy+EmtXwKDTrDr8LLCXy9Jwp//guuX2OFqTOnNCIrYWFJvojl
nGTdxglFlqoRL5/WJowl+zwun0bJip6v60eV2zMYRd5N8TXDCy8LYo8Aaqe3RTPo
NywfwZcKDXQ0mzkTTxKY11f+QJHbuVttmugdx8dTwkMNBjxlG4NzJuIsLiPVkVmA
9evZvU22sCr/suqfLYVS31WqrtXB63s7NtTXWvBEJQjYx85ylf4KdfevWnao4wx4
oGKeF5KbBUvPuK+Siw28Gjh+x6cewMV69X3Z8jqK0YsJt44afvEUDyaipqdk1GCw
SqeE1FzS9j+5PBLYHpuddGSntZURmCbHF0MPOfSGnkYkXU1CvNxvotcyKBjZFlIY
I1jIzjC+hePAT30BZd2BQH3BC19cEZWTfDALTmcNFVIaIpXcVX+9eRmb+GKRPtS4
iPaoxrnMI5jgwpXEGdm5lFJvW0/xFKN7p5HpyZIs6CsWbRSFl5+fIHetJsdkJV20
xwrL9f6ldzkezOMMt+iNclbgdHiP75P4N6/SYUjAJvXxL/9r8tRWPLXPZ9s20XuE
8xoZzXDftjKlZ+NUSySjhnWVAqhSqRuS5613HP0ckFiLI9mXspPqJpj4LRtQe8uR
2dORqkuGRsPUn+NtrB0mqo9Qez3dnQ7b5eZr2/Ob2ghi/BuKtVTbTIk2w/9ta97y
gUeR/HKbsWiVca0nXHHzpF/vjTIpcyrSxvqjqc5jsRcHeB6S39Ndqa7EuNz7BBF4
H8K0d976VmapVgfCHglnGKSeBsjBc3t64EwN+yI5R1MiNj5bjmYteeTIHR/Kzhsw
Wdv/psBOAcaFJHVSm560O3gsgF62EJaPhZ0P52pjFRRv9Bmw3LJqbqMUoPr553Sb
DC+aPgqPXG9+w3oOWjAPb5WF41g88WQb4qoGGngPwSKI7729GVs6i9IGXt1/gRpG
vBF/xmnoKU/JxC+pSAU9j2wA0/nfaPAhgO4VtA/kSWobfB8Td9YWvTLsBG9h5AM+
NW83ppeR95NfHKdp9BmMp+bkst3ekp8kBAIoq3GljnQtj4sTGiQsBlO84Ukn77HD
yNQtvXc00vxspnOMa09KQD0gaEuvLM+vvd4KnsJD4kThnEzu+/pNYhCgrhyMdwzX
FcvAG8glpOEBinqi69JPSAESE/WxoZoEajXD0WwjjW6o54PtUAe/11yet/iszLcD
vByanf2eepP+Xp9n8W+ODWn9ZkQvtwMU6tuD6JYK7/GRCPEp11ZEbR1rWClZwtrl
v5hiDkzk7/UD020EOkHIB6KWPt6PSQPU/9qvibSchoXUGqFIcASfdfvHxUpfkmYi
eC5OJBbeV9uDdVLRTk9uSRzscbBMx+bon6ZNUMZQFDZxbWBgZzM6Na+X3ORSiGki
n5SDKfDfRcA2nQ3ZTrKD0X/lTfebcu6PeDeibrkZMtozMQTXlM1PecMrhsVXKYvd
gjPlrFNI1FMXfuFVH0FZ1Lf/Vy8l8cHD6VUX8hpRTnMkQ9z9FMp22VgsuXw/8dfA
yImQxPpDTYZPDdCPLcLnoQ5l9VIrrwa1saD2PcDeBz0VMd9DdfllTERUvBwXss0j
3ZA4dSg6KPZpWARtThyS0geF79jrDrFqsiYtYqXKjiWgun4cN5MKufpOPAi4WXOf
OKgktES9myH9xhixdUBgJAbF4ckGQXaMW8j8tw+9anAxzMls6wYfVBhddrxnjGru
J5z7qElMJnWdljN1v6ytBka0uBgeLW6b+cDwU63pbqnGsPo3ZGnBds8EzH59XhKi
8D+aButaf1rCd0xb1nxuj0y8XKiXY6DWbIM8qC7ncC5A1TLTviFqLS/OmJMJ//Wd
HjvFUWIy1UdI1cjxN0QBuptAPhjSayOfA5a84j6aiGz4cOTTcC9lDPtNZBaqxorD
d33zCyMUJ2ZWKTsqPpv/dCP7+maXSP6BqAHX5Cv8dPTxuNPoJKX3n8eqPFmelqmZ
P+mvDQlNZI9fmJMaEvh/if1qYaM/uH63KtGlIAYpH7MZtmX68fJ8kz6+x/q98YXQ
RSxMkXiqt3RYGOz9uv+qKHOLE5GCScTjex8bIk91EuJKhbMTakZdba7U/hZwwBs3
/VXyraVxUm3XuRWgd56j1WuERW49RWjy09/q3Rhsuhwi2EgX1CTW2ZEWor3gdxVf
i6NtHKCkK4KMpV3oXcA+cKC0Nb3n/PS9qLeRxDUEST7bIpbaATQM5nO2M9YKGfGG
1wIJDiIoNqHatHJJz/kOjqTlyG9jIANSvWWIO2GnnZqYmViKu6aV9AIGtcqg9sgO
8n3/yB9XhFll3D+reaTxHLuW+aqQXZlckYAxhwU+t70Qhx/1keantnXu1nnXgkIX
mSqV19+SK75eLTq4ckqFB1tTbx8wgQjoj1HvHo+k9Wga0qDnUMLO7RDWQaTtZeeu
JvP9qoK4K6n6hxjApuWJe2veItULjDfEtqNmhpHq0AgaL6TxWs/YSQl1RdWkR8Z0
io3fL7PsCir19vp+LO+zVQURRwYGAj0ND0jrs01C/94e49XYri2+IrBcGmVkZ9YV
Ys46K2nuVVSQI5ieZmL3DpmxlXOLoO0EdZ1ENq0iSAnRmN0vxRU6JYrpXLADQS/V
0MFN/JBZjrZm0OblfD21qz+GUR8Z+CrUwFxYnnDm+SovjiHl2Wlf7BElTrAI7l0t
djU054COkEKtG8OY67aS0SFSwza766Py8C+FQraclkRc9Z3VZL7yIC0gXgh3tOS4
/2Ag2tJV+jRfnfeUSJC8LdT8dZZ3kdCzSr61QCxTsGmgFp4cnOfmJ7ekmVHueZAI
Dg0OVyYGhwZu7mZePSbAWatPIFf7KGeWG6kFQVAnrtZfTOWeWj4RIQUiqiL328WX
7yOCM8vzxotnOZusjsx2QoONxLptLiboMPTy0BCy2cQxlKogUEOGzaLP/sI36TxB
7y+EyT7tqtOnoe6FITFp/f41fFMSumFJHB2RBJ5QxrXo1DvBtUEnMf7tKsp9o7fU
1O/Nx9mwAre6o9I6c2KRoE8UdaN2QE/cMRDrWppH+yhPHghQHK7HFPHOwgV4qTcE
RSDUl+GpUAj3L11UK5Y58BmgJfF/WtWQZREVj4edrzszUt6yRSo4Hky0AmK3GyoR
26Kj60TPCUjLRJKCRcZ2xxXEeNJyVYLUzCLwq4vS12qPzeCAMTDWDXt1wx0Gs80B
/a2NhLo/aIoGNOBs3aWS9DQ643JKxLMFpxk9a880mz1JjOyrqwODZeatBFo+mF/f
Qac8+olItshNfY4/FV+vv9bcvcdnrtxD2pDGHoWM15iblMrm3BnpV2N43GqnZGej
xQybpdfz/kIsEwZ6BgEyS1AVvT4z8KwAgF6wf+Hmlpanf1DdlOxtN4UlKhEryPwy
nC0akyMPAZRGwMSZ7IzYJeejdrojRHvREdU/toxO3StTetSLqaLx2vFVXwL3/kgT
O3K8eynsgA+N61vYQFrYh3vjjh6yFUf9VkLG8Xkrb4CwlAbaKBcCTFZuHCPufxma
eKWMQYTe6MGaXQknys69jeGejqi6YqvGqLjSHjc7v+k4RLlnA5UNv9+LxLtoHmhb
LAdQzfxCD1Ep/gaXgWbVoC4afG8ed2/Lf9okFQ2U0b5OTcJSWriM8HOgife2wN86
g6TZ71JXAZAqmWPIAAmVWyO3NeK7IQp3eEAEhaADqGHxMYKGjW6rh3Rq4wDw56nV
13pr0tfjkKqVmKDS/eXJbYMfu5LCAYnmXUCqjZtLgSNXo11gclZwpF60wQt0Sx+g
HHv7Jn4ctFrQENsaSEOKm8DGgp3nOrDH5o8a7YDyBi7Y20HqfzR5cQbmb8S+qA4C
BDzU9afdKh4daicWS3oXYTq7jSeJhTUxRw/cfH+WCmuUXOP4Cvy1rqUY/8Ay2DzQ
A/GqIZcdWWuwYJ5VhH7BRxjOI5PV0wHMHv53a2WNKReuok5MhzgQPiwFHnK8Zy7X
la5qI1WYwoxg7UlmDiVb1GeDa4MwSXWpG+3Rj2KjbkMG+SKv0FbauOZPCjTfGvBZ
Ci7An88pQ9AC5/zV3BaKiXzXBnT9mz/1Tm/GKSlNo120PSJdyI2gCBkpHnxj9fEp
dtupwKsWtfLooL5mZSJPzLp/03L35oV/uX4z31mQcRmGlndsS3wcF1QaeNICUHrx
PeVjSNM+o7TdTdt8k/IrMQA/2Sr4jXMIM4FCVQcouzfKvRdRh4GRyemW1mQ6n78t
SshAEJhYvMMNDbYTj6FE6GyWdjoNtBXLfOjWBAq+4dsY1JIp9GWGhYxGoxacc1eJ
XOAuj11iMeDb/DPOqGfTy3g1foq+dzz19rBZDnUX/fbovEM3XKBke9EhHhtiYN7f
l2t5V+hgdsPT9KQaIIPqAwcjsbLBWoRbvuK1zRdmw0fzNpl9sWi3evlBKaNm9rzM
DVQG7dBeIFjFaqN08KYf85vET6opzzA9fwB1S8+kfBO90wig/q/v/HLPUqaiBzBg
KmWwBpt1mXI+ZmncrLKabr1MGj4cHhkKWazylAywnsbMc2FqeheQfQQEh4HHlbb1
z3y3kjshSziUAfL/Yr/tDlMz4gggpZs0vjb04a2UvPM6NyV00+qCZjCF/WT9Z71u
AeIail6veiMVXfe1zQH2MtD23JZuFeaQ7eDModDbdhFlkdCcbIjLVAvS8sMZdzTc
/6rlXNA1HAxYcnq7Z7lgoUYK46hc0nobKfQZPZzaHl5Wm4eCfs70bhdjbiuUzAxV
LVKttr24dg/z697Z9erUnr/vswax847DJgD5IS5yikvyMilcDWEARGq61Qr0Rij3
YM5yvDo65OhbqCdMrCRf0Q9dNUbVv/vT25LyDIRXqu06yNCAIFjeb6jA5MiHxDN6
6fcCe55qor5ZFHEPAiFBNPCteS3EToh8WPaJ6lu+bToSuvOpu/lS9ak9geUKDw0Q
Kn2fKrLdlxaO6zqN87Xy7vjLLoodPkHsEOoU4QMyCOk5G3PtuGisN+6TfUr+4ZK/
9/rLaF4z1OBazDhYPiTUIK2PdVRpWrUmeGMPpf9Vm7Q6CXYJvF5aDOLAc/NmKH4N
+NlT2mxm2/91eiMA1I9J8xnKMgkiLC6ja/0agDk/7hU52Sr8+eWSA0feOn2kFm4a
OXe/VQNNm+Ap47tgYSgx+PRbXW6UEbb6wBKvOehqoTRcVsaCLMffmX8YbGpf6o7F
9oVVuDyGlAbD6pCpNiro1RONxztL4+q3p3JhDDn/Cn21iq7KM1A/83ky1bI8OPQR
fKumW7Thj+BLDYgyU0hMZxWgNjoZ1otXWzwqCG1haJCsUfGb2YN7ZdK7eOBrGqrJ
STA7TONfIJgA21zmgAnW1vTVOyBdlU38ABpg0NIUPLEtiWB3cYipoIVEkMHJLMGn
/P7swMMzZn03Lg+QHrh+mpKuaaM55Lm/kJUG0TqX6VUwvF8qKTczpuN/MPS0hqoK
5ZfEjTAtEjMkSiwEnUKSzQY2k7nqYtNQVUhKrO8L32UB6xOD8tVIqHe7W8WG3l71
apAL4OdTVvLAs0r7ulosKE6n4qAeqxM4mfw1cf54gjMKkUz3SUqUzXZQlApAW4eP
z4UcJZYFkiPIo84Pyqv/DLmNW7/L7dni+orowsxh3Rh8VZqkaUlngB9qOYieN/bt
FqlwI+8Uc/xy/O3Q5wVcwLxq8pibrzRnxCBJNC5JlGDZN8H5U3r/7plwn76LFXst
GhsrLD80s3cVnEWI+8nX/5rssc4XDT6WX7G2UbRwrfDFSPXTFDA7Mhp8nqKCGXJq
Zm4nm5DL8yes79GYYT6AM0DY7RVLwHZ26DGe7dlKIPnuU7NvcOCytrRwfbT7jO8t
Admnocr5pgb2bSyVQiBx3l1dTUSgMXhkVuk1RxLgmTzz12jYXsyj3URPielehtu2
3MoXuuYxoRLK9XyFvP4St6wboGWg9GC1ej8S2zrUbWyznKNaoifnKfuL2nroMbmG
f4y9W2V9nOYK3gaS5SKDPlruMhadK82sMG7iMT88kNovsJq7pwaFYFpx9gJPlXIF
fcrozKYDYtfMn5G1F3kPE1xmUlAc/aNRlqb1CAy17651LToGMKjRIFcI1X65bd6u
50TXPDs9QC3IDWjP7PwInC9LwSGd5xK8XF3NqalhEbrg+2FSg1CtR9uBPXr3y7Sw
csK768JkF+nf1+kJRlSC8WP9Yz5GJhl9v+GCkrB7jAZFUMac7dIuAeaLBOop0YRy
jmYL+5cj5TwVB2DX2TIduOZEjKojDd1/D4xvJ9QVDxdTA8G1v4IPKZC8JlTIDZBR
+jDhDEGCJRyFiA2cCPDgSJHTfNNkuOkQr+yTw5uWrtYMAOVKEKE2jo1RqQjCdyZ9
709Hde3hs5cJCXpsjOcqRoKRMnIDWgN2H3TyK5r1j0NmD0su8Jpf5MSQrReREhof
2gVlEfUBLfW7g5NNNDjVFvTv9mCsqfBszHzpXUpqXStJl32zGLe3ibAJfBJ8GSoG
f1ozcm0FWNzOWAkiRH2j54abh+q9So0R1+w/jrY+nnWy6j8Z6pevftlleYVwseoF
ujunN7SixfKwTcFKVfz9zTaI6FvmPZs4lV8t+mvFmnfzoQ2pxudu7HbbtGXhc668
SmwVbdaOibTuj8hvFzq/B9aqMys8DOwmcVuWGD98KCUscT13XaODHeAGk8bWc8bd
6YEpkLahRY3Oe9m0XeBHU7jpwFXg+mbHkvPZMI7WrhFbpCeSpQP5iQoYR07YmrTw
R5BMg9xhiY7zO9sA8sdOhBdMJREJtXm7Qg8KIDopfZ63y5WNGxSqqokAD5YY6Q0l
jfM/XgMX+nNsAX8PVMA5jRVrRBt+o7hkHPLr/3bi8/Lc+caUqGVCZTZUWmAyOLVp
3WCEQGwzwSVjjp48lurXz+xyl97VR+swuuU6IiQevapTgz4S9ztkDvENB8syTBoZ
9Pm6tA2IuwuFTxqC+/qJUUHZx7IrFDOuVv4sWD/5qEe2ODEF5cqjd2LoUVE71SN6
STUKXY2mJm4ZR/utAjoZ13UD16ah5tVu7w/YUaO9KWkX7kdYPv01EsXuyIT3HHE/
JeGeomr7Pq2NYeA9KHzYpJLlLlgwZaAImzz8Fpyu2f8jJlbr4rFWI14PSAeguSNQ
sOszQD4LW6Sq3Pc2rxOG7uR6SXvh2Qg5eL7i2c3onymwwf56bZUmi0Tc8MBazkzX
AbvCnRG3d3sM887iJo/Z1bcgwObhMCZZVIWQg8CVWJ9WaU7twiXp3bI7wRiw4P+o
ohCErJNk9O3v+Odq9djQhAZSZFqR0vw/u1/iRlN/nx/r2egdO8UTgY/p/2KQQKcV
5QqeVV6yp99N8lx6Omjo5q++89rLqith0pM9Ogmu1Qead9euKHBci5DcliurRXVi
dlLzzT5uK2jeVrgtAlrHo4zIHkRZG15vypEzVsCiCLvYCb0iZlHkf5/Hzmb3Z8Tv
hr09j6+mnHCiMaDvCl/3kzxIy32D9dOYa6OeuOclRZnc3Wsqu25+kFkqMqpICt7/
XY63iVJNTmMZREftd2C7jWFrVZ+5iGJ4SzaU1Cq0aFMxKULlbzCxgtrOO+bBTO9E
gp+UWvSKm0Y4HTL/dj0V2440XECGmLaGdP0/18t7fgNQhEaCZIjoZrqUnI9p32Nc
qf1Q3O5FVK8kycQXsW/p4QvqZyKUU0wz7EX0znAGTFSyFVF8NvR+rTXEB2z5hIff
/slaiOZ+tEgdj5tKEfgnSlBHhMmtMUpgT7Xhb1DLSWgLrXaHhnIraYlp5DBQS//I
Jyx/qSSqY9TnZQ40ZOWgJwnfBorIx79HBundtkbPmlfBJ4ukJnSjzz+I8SPB5vvt
ftMXSttpopwdZpTV3nUsfPrNcnK1t2kUNS4GFD5edRkwWKwzCejunBYGeiWruE03
BImthCKEsB3sxELLxs2sLzPC0u+AnLsRb9XxkOb9aYlVyeOFP9obUy9EKM0AsOwh
GypzGf7VoBGZCKuyImatftY2EgfjLYZmqpnY7y81yTPgYtBvMB1H6tZT5AQkFN83
yGHKCAvytAhMoA2HZErmaGjDj15kszvSvIry/QKRYpcYx3MjrQaRzb24D8NfjCpA
eIn4zfSOhnkFSX1gsAzVovhMTKFhvJo3qlcbLZGtSn7nnQYFIs6KuIPXh3T7nCbN
NiXuOioBQBeWMrSklFHupkS0t8lS4UaK5nkLB+u4WkPSdMGWSuq2Eab44qzgHZ2Y
beSf0RgOEK8Vw/samI71oSlkOkA2YWFlwZYBq02JE8XKcI0QmzBrlo5a1BTtkC9+
hHvpvFKpYKYUeBY+3CzHWfN57CL+4SpHG3U0FBI1PJSKD6Fm3RngA4itVU88SCSD
NIL3BhlCFnyInYIdq32uv+l3bu+8rS1Dua+cOposf9X3cvxArSZPZg1vs6kQCGg7
oCrfh4e643w5FjtxVJf6uyWkh7c7hTuJNUDuLcujbu8rdknRfhDCMGoyBAqRWsfR
clqYscBzpBb38kO+LlTV6TQUOo/+2UsIf427RVKk+LF0nUdEI1xXiE1I39o8BET3
og1rNfeaKoU7rQb4B764S8TJ6heiHj1x0HrJENhcCjx8RUAP+RRKSNSDVBY9QDmG
z5Ow629VSwMMdH1ebmATtHA8E4yas/pIePWOvpq/TdWdc+/6N6g6T4AsIapUGdTI
IbZUiWOYGlO11Dd+vCwGy8pblMuDppynMtmezH3pWFgFFVG3YnMph3gfc+psbcqM
DA41TozC6CaKTnGuYJzfref4U6krw/O/wn+6uMA34EpH394T0XCGisI5cR6qAZXi
PtTM789iPOp/+IanVP8hzqgLVv9iXJudD2LxtrAa4lpYNIrzCLa2iKB/4uccCyXX
4gRVJGeNRsC3xBJuUqjrjLijgv/sCuiwyASMMKb638y2je4WCT870UxdH9Ck2LDD
riOSFT6mQ3aCCPOjqj0YIPOTMcBEP1pl3dhqMeW+PVP5TXfMNNL6aRsKkRi28fLr
g1yP59vl9Fm7xi88EjSHobjS1MXchZi6TncrzZebJUV0eGwANm3rfloNDYTzD/q7
0N2RFQulbHZqevDmBSZRm0BZ5IV24wo0Xm0PEyAQeEHO63Po7xeuaEvxoG58ZVna
Uxf5TI+PZOY+no8yHRUWD+q8c0/ukubILqhds5GAH+2Cmk3qcO1iaUB9JXENSCep
IjXoH8SpyHBGT1iOtKcaU6HbK63AvUFnkVzHt9WB6g3f2Uf2KJE1wmcGwY5IsyZU
hqUddSufQoh0emzsh2wCQMrQXX+uQxrZgJNvwHTWcVPqAS/VLQrjuqCj+bVeL2m6
gfmXOJLwXbOXF3P9V7GczIraMosrUiPo6MBjGXerlGerHSzjghNSXjrb3UJkuv5n
yP6UKi482CJ3Gc23BYyxARKf79nSjChbfeeaY9y54AIdAgRf9COv38fR8dai3oLQ
KynGOzbrTYCB1E+bwTakW9SaAVlwSyw8MJqTl/cq3YdP5zDidTw395tC9zZXWEeP
g9ET6f2bPawwzWnERa5gbX+EwBij3+1CDJzTm9GUaF3GEjb1NcT7Z1L/DXLlFM0T
EKhpx8ExR1jZGwuivUUh147AftntZ2F8LiRSt7iwpDhcYozU1ilR7wIOyrzOxXwS
Fj8Xmko7G88BwMmMjqmVYnFW2BSIvX3BCNeQaHeRxuC5tNvQRhTkfPj58ijwRB8V
ykunoE1vfnGRbI+4Y6rklQ6hxqDkz5Eeegqy/3QPMT7bc6F5wfbcE1H5MNvseSjT
egPxS20WFwbjwIF+7Z8q1n0NHYjjkDElLYjuNn8n8HvUrdOaA93YU2YSq2a5HuJb
kvM7in4UrOd4bj/mPsYivpxJcJtu/mGO1uTy8qrJjC90WeomgW6AH1v4yA13o68l
fzFHeoLOCS2BzkmkF4icIl/mfgB75gwYnwYhjYfTLmI7cbNWoRQsmaqhxTJSdsvL
6pF3Sx0rvK8bQxusk1Snp/0RzIJGiEV47qpUjXHaRWrc7QhAuhT2AnP1G4wOSnRV
Sc0OyQ1oL4LJf5kCKFArBH6E7c3m0TNPuciIEDqvLY+Upmyx4iCx27/euVjuTZZ1
DM2t4YEdYOmG3wP4/EDaxdhpE2Cs4LkYh6qYA3DQw5WSUlqWMlTOzFgxW0WJbe0S
O5liuxZk9E0LCAUv8hNAaYXLWXxCru8GD1AL+BlHH64y6CvxnpupgS4gpNV/eiHD
p6Ivmx/+NxdjKkAyR5yAsFKRbZPFOASEhnHlHXknJ9MaRSigKkv73bOpLpp34QSV
Gkocw1XLhYWR1HrHYBgGevgJR8whpT906c/CBzJPNwFiTJ7UXs3RUQqI3k+fTrC2
u4XDVri5q1xch8nMuckp3bE1Uro1+eyUBPl8gsyYh72lYTKCoylyYE0Plyj+NiGb
zQ41izohjKUkSB2sf8HuwBo9gTlZZ72LR+oZo/gHMUXlWqG0tBffHxYOazxmMF9c
Ds7ZpU/bafPRGd4GPDN0L3iRGrMLf2fObidaV0Ndev+CB4xWTW1jZxGvs83TxniF
oLcdAQwjShUIJ0E1G/aDYuMxoCOYOjWrYTJIOidsHATn/QfaU9+ijZaellpe3Cj1
Ih2b3dEerE+qA9nP6s1ncW2p6MuM/9i1VJDl3Ap/tGTw8KZGD+LAsfX6NSIwp5HA
eSiRyECd7RcJImH3pdRiZ1B6Krqx+TFgV/KRZdOnuFi+HZR5wkU1KWC6kb833s4D
xvh8neFTvHmy83N+EQwq1FxTWB+p80fgNheAwFzsyiSV7jH/KkQ4s0l3OzIw5xwK
3oeuj4sE+sonyJY6LBUW1HN2JYbilUtfkthkRXE4t7YdGoWVzHbBIcYqmj426z8F
gdnPRwl3dwLwKn55Ctf/IHn//dMNmJP3gbfn2rApff4zodReejCZ1UucmXssCCpi
RaUV0WgYsdK5UH+3kcMH2bJdjJmAqlbIIy3KKCg/iKf8VIVE0bwJUulsjy5TV93I
Ipz+8F7TERGVJgscoXq164nqMT+HCLZfVYk8roSqmqE/mtBCY0CXJL362s1mJdPO
9ep34JouH7e9WGHyAr9iNfnrqELtH9phoyVRGZ4IxfPjd/I9mkpA/hSptKXg+4ta
gUq4AT8uKOUYJGmM9gp70rISFxDjOLrIncABpyQa2x758yduFohdYnPQMMdWZ9I2
FGv6u9NS7D8c52NOLrAVj6FKzClHDME4h8IH7cjxJoDdb4lIa7HKS44dsROJmpXY
MYJkGl5qJ0NeNgLOIzrAS7Cd1LmyjLUFAXN/SLoPBiPkluhnuTsyw7mdCZyDqh0t
2P3rHUBCjZwfjXuPEWxE2UgUluROSi6Xb1n+dWqXnGCLpTkHjaQNZpei05rkFjh0
YRJhPAUxi7MijIxwLySz6UwQfLM9h/sQIAn1tXqNm3iE0R2mePKaXlr2oWBTP+De
KZvz9h9tV7QBzWb1q0ZJA19BDGXKH6VCrMJlCm/60cS07X+ApGV257vc7WZ25WiA
ZT8qZ6VyU+Ze7hx5CBiaPUmrXAe+m137Kv37IKj1J5LZw693r6rOSb9AJUboEY7F
fudb3mcvsSu9QibEDaXGGQGZPffTtELFBc6wzu0YFQTT3E1r0lJq1vnid3Ut8po8
2iVlQb3CAELUUSeCPO5ZekG9IoLym1tEW+RxgiS5fUBh9OlQJGey2C4Gh1O1O+D1
0GLU43gXYewgHpV2yKH9eeAFUcMoUxsQXfXg1sJmdxPY+Zz1TjTgPkhDR/Np2fk5
yWtZyvFsqb53szkvPN7W0irA3hplcRBelyHhs64hXdVxV/ocU7YWW+GoBloCw/62
Ckt9x/wX/0vY+p14fPKzORyO/OxacongvMWrWPSh69qvgJ3JC4uEdHq6Vz4cH8GU
Qp2LiWDxsGzWP+aMKI7HXt6w6ezm9kIPcPwP56qjjHjdlzcCOj4LId4VmMofnvXd
15AZ2Dj8KFWVwhELJBEsSYWOHgts0c3wygF/HhihVPpVDj2wwOauc7oWtttzFyXJ
gertynyqIktj7H2rRUnRVt5rqmlL45P1S5eQeCz0HyxGBPMu3xAFr+gkrL6aZJEV
1kyG4re3TX0YBtIunU/ZAX2VyO2ZsQkBDwkBpcpnayld3pVWXf7VdBVABK5TquL7
exNAVDng0C9JLeRODBpjTLESkMNQ5Xncseu/1nIY+6czSK5LV/5c++VvweD3HJtV
fc76WyhqdCJK09vbB6GehGntpu8aBqjxW2LS7MZGX6uLySVeK2fIqvl0Uj18qg5k
v1o3BI5fqXs1bWMcAf0j+JaJTnFH2Cax7tSnJTFKSTms1J0ArIW5bpXpAFF3sBpw
5q4Ur8vsYFNcD7GawNIPRftLiLlaKpvviKsSEGHtxLZx5sV/lgf8zNNyNBS7zmTX
NsKfeIyBJQMiLrbWfC9juv+S9F+HSkZtu7V+k2ai5VIhWlvY3RXKeHOvfLPamXXF
6AF52dvdxZwWUq9m8AUjXc9dSEc4NACjz4fvYLgIjYtTGLRahHAkhNM9bYowvW4y
PcRvS0eJ8UdlawiHCrtHOClUK8qQmyTtkKblGqR0T0L/B3KWk1MMQGsFHQKsjrhN
plzLsxBdx/kEwJAhvcMBE3NTkw1uXKKzG7aqmTpojugjaYRltNjicB6DSFieIjj4
h6+9HnwBKyx5yPLeiSo+KoCjgvA2D9nhKeW8dbZIA2zVUcEdfNIXeVWaQExAjS7S
IaRhaaLz14gat8DAXr7qIez3wJZcXEf2cCPJg9K/39tZURNj81u9+65OTaAGOvCT
oQRe4TTEkR6kCYFXil/rNTBJehiX7CD5cGAj2ON981zCFb7cLSDTjScC0zHhE5Ft
dQWx7C2epBiljHWv5b2M8zFc1MvUi+Ys2+V54/PGdHsYrdG8jZc6NH6/Tq25UndC
yr73d/VirBL3IcfQr1VIO+eU7Go2/ZfWRqd7z5KZOM4UvToTMEgGHI5+Q+6OprnT
qFBMz2pCKgs0n/4DrA5k/JiWpCOzyH/zVSbXmf8jWc2EY3z7wqelSXbLkPMVU1Sb
84ewAlgF95IFdxDu6WCjLSvo5Ir8r9pE6izSEOpd3m32snPowP2glrU9kJww5SRn
TeXgWsayocM1ROOne+i9EsUwR3ByYRqDvCh7p16/dNC2ro4iX3NJ48f1RYwOVKvQ
iejmof9rLkZHtzwCH/X0oRkzADPSRhQZhN8B3K5zKDOP/gs+j0rJkkaVj3C2MIqY
0BlFDaSqql6wY5hRcK+WKLrt7X3HyUuMXsc2YxRqr1iSdb6irb/ogCCe1f92DhMy
CNXBYDrrBaRwBif+8Wnf71I2yC50l4LrCbFY1kdPRgiVLNN5/meK7f7/68uB/6K5
Vsveyz5H8aQLk9PgS14aeYId7E4SSL1vfrYE5Abn48WRpymqIysj+pvgtNg3iCtp
W+qyhTt9p7OdrlL7Xn/iAavwhTuSEbw/+CXCIPjphj5yS69KAlh0X0GOFWgkY5az
zi77qWMxoetP/OQLGxwMHrJpdYOAdqSre5ft3eDmSpd9xII0ZVYBlkaa5BZtGUDh
UXjFksPBz4ZAkvYze7QmrWtUambyZvSTObMd4uOyaLQxLxCf1P056CZOLDZN4QEx
n3Cc1dGlzVWqzZsW5UDfjwnX/I0v51n7ZW9NIfRfwJfqX3vcHXRjYhI2s3T3s0XK
K+GbA6RpZtG6x/tX5mUe2uS5euYQVBMvnlE3096RunbZ26gMMrx6UmKjFlOv6ouo
C7rRb8xH5l+KAzeszT2FOPx9jwhAg5gdjAcNjsvD+0+Z7hexOWT7EOUhixkah2Vl
yCZEXfA/2DZt8eLjKiCFm8GYsuf/t8qEkmuw9DXnSEtLWBKk6tfq65E2lISFBKWp
T0Ok11XBhW/dACIQNVSPjf2mciHr0GTS+O9c74xGALm5fjjnQ3WiXrPkK9eEqDv2
r0PZPXbSlLFsvE5cDWLOl+bS20x7s4jyvx9nH9kGJN1qGHiooftLvYn/atjd2AaJ
cFT1Bu5oZelG4oUcOR3WTzOuHb4vgkrK145hJofSEe3jQ/Hx8u3r7dIG0DqMImlV
NlSlHPSg5lpqcQDtzWOsWSejCrPAxBPl+V75knC90NGwtKw8PxlEpNKO56S16+jT
85m8K/1jlZG9EwrmB2R+gc3R+2zSKZQZsm87IJJzv0sAXO3mF0EZeIwPwFIZ5tzk
472445sZI+BEtWP4eiC54LnqUt/vtGC7Bt1eQUhei0ll2tfY0G8J/nfpvjar6tTq
iIW7HUjz/PuvGDUOOamHJpuaZVoIpgwoLp0JuR0Rc04bKiRUgDcJ5pBoHYbJI3RJ
lwjEUFouOjpdZHuY1Vx6YCd3nwtGEX84b44SwCVKYdqeDiGKFzA2K4LlffU9TMff
5GGDObLzz8yXZJNAPPnTZpr81k6+tVg7j6RIHW5Ztpvuba/yF9dtSjvQlOKZda+Z
xOYPebMV05xsExuVNcOraLLwey1RoTK2/Hz+4Pbg1JVGlBw9gWoLIO/4KS+6niur
Yej0t9tMxi3/ZpAhK6K8yerrDLCYJs2ZEzisvuc+kSnYGR7SYAKtUnJegttMA6Qk
J0A02I6smmyvknvHVd60wNJ4HYZWkKq4YTGNZynTnOB4exiEcCxf2ll98Ch9zbjo
fOKsRDlogJiTsHvCwxuEqud/+WVXLGpy3Pomvky1nj0Jb42VGCCZ0bQz1CnfQ6Us
0A3RZR7ixYLfmq1NSVRs5/w+HXugj7dwDkLSVf43bxG7p+/0lybqpo9BLoxYhXmw
SHU4bbHWVz8J1T7f/+5rNN+tXQ+RG9N5h1KjMtpFq91w0eExmW0/fYWLNTteNfbx
Y8mV27pYVnulZbc3i5+PdZ9ZRQ8pVOIHzlo7w1jCcrVi9KNc68dP64CjmzmS1wXy
OspSBM85F+AvCMETvGMl9TXwYiShC8cUb4r5wT1v42BRMlqC1+3Cid6w+Swz/2wg
D30p0bgzJLs3br8xSJUKExjiwL8s/w+LKP+WH9pGp/k+kw18YNijyg2ZnxsHI4GW
5EfqL9U0pRIkUmZ5lHTYMfmkaaJi9dToxTJE+8xLvFG5TKCUlKySE6nE8OzqG1OC
q3cr9f/76kL0DxDXPIYjA8RcE1sCcZjTclU9ntJ+XC2H36ScNhn1v+lxCr2Krwki
O7P8yDpmE2c/LGcDKKUxluG+MHrj7mda1fa81nn0P3qL7+0MMy57TA54psri0Yu8
Wu08bPFga4thgRhdNAcQfmtTgGiL7p8QBYWXbVPsDU52FBulCHeiQpTp+LRuODt4
k/3ZxdW0xQZS4rfGkv7FtwSOV51Iml9hfFGFQ1WkEe+NCbbAy8Pka0sOyNLXYMSu
KviDPHEbA8iTIf1VcVKJT2ht8RS7LxEeCCIcZkBPdPVMUNt1iN4S7Yrxbww8D060
UyR1ywKsXfj9KuR6rBkR7m22UMlrbZ41j7c5oSrd54yPfkpqX6oM06VyIfK/jYON
iSDj1kaw9eti7jfUcvDPDke0qAiAMiJjCP0OtNISFBV8sQq26YCEz/6yoNyBx/uZ
MJo69Wzu91VcvZqRdBC7p/Ll1QQsVIyfzZdzbAUKIOlO7itvJYDzDUsGW2oxa89l
TD0Fme58M31xna8Vpn5zybm/jmi1+BD0McOFB7Fkh7Mf4/GKj2YV1E4PVO6ssxoy
uJ/Few7JV084TK5dVMeTvDKT6O5d26Ypop2T5n/TIyjXCVAV9qMmveRiq/A7YRmg
unMzCE2fd+eIuIR5JuPnyRIdItsG5gUJezcCFY46kAqvRq39Qt5ANjRgbUVH2vQP
DFNMpUd0AisRk+x77Y712wZ5daWBOX3cNL3E+6QrzjYjX6Eg7Y2EYBpiCOJWL/OM
au6pVMZsyc5ivdIep8n9hqkYqOtJzqNLBjF3SvcwBkJbxzE142THOcYJ6TD3NNbi
Oe1w7CUUCMJRFu+JycgkjhkQQd5hxqpaM8tqtD/oFywV7xyUGfxYPEHpdmhmyGaX
Ao3vSJzYChWsKMnv5HB9oGPrBx6uVvMeSXRhY9sc3FiDZ7JT7bWfsPFxUd6DQgVz
V+adMsY0iuk3bptdjxHuFEHvr4PhYvHr/iYOW3pBCDK4/J4psWpLNB9YnLukzzkQ
2s4BVkYoGaJr/jf8nzUlvFtLHl+Jom30xTY2/qp5lnrRTU/+0Gl1I8YZ27VIkoFh
O4snEhfVrEXj51wdPsW8Baw0VN6oD4ckLykxTJzdNY5hAnUHqVZAEPI+miviquIm
auU/M7IIrzLD1VHGqZRY4Aj5eWHYbWR0GGAlEmkHgf2h470KseUO3QCMVkeW7oie
Ozeiu4YUJJnw5K9jh+FsJmkX6A0/UKmfgqFV2UrPwrOQLpv7CumIeHTx6Scyh9Gn
mZgqI3+UvN7ThM+gmZiFbKCetfn9p3AS0Po0iUwL2OHtXFZQjaB69qDKxAYRNK9B
V2bbzCeT+1DZfLZzQyoTV2tbC1sBZBkNkGVUK6MzwIvMmCto6MQZsG9ELpekJgTl
wPYJTKecPwbA+CnrW/svflxj6L6WH5N6ML+i2WpWdDpZsmYQfUsLhBVjqiv8G9Pa
FLN7qG/Z4hQ6JzlLhuSTQRgVEmKDtKCKp32jC0pitvAfqGXtVtz3fPpIsrTO6lVi
Xt8trAYBsUe9WGFJ4cs3QaFxMZlJ/ZDuaRkOqyuu/yl4gVmBO1qU1tKjmVAf/z6H
Afnph7YUMB6SFpF/VtrfAsvxo10QuJtfiTy3jBb9tXTmJRnsUTpbn3VKw3qdShjm
0dK/7QCNMjXyaBOjWentx4T0i0JaIQcx7BirenLz3OwOErX5pMggOKHflAHIy524
Rb5LVnbDO06v6L/e7ie0YTXQ2MNaSW5sSAQtcL1qp0NDCXPFOs9FUHk06WZHfQbs
U+gRIPSY0ssmgcBceikxlfL8zipiCl0ETiL9mvQqAMnABmRBki6rKdJ0ETuI9Q9L
tzdQEBvH2gfHuxJkOQUmk12pCKxLDAszF9jA6JueW8yJQ7t7nq5AFYJ0X190MQI9
oKDqJvG37pMt66uSjBBksNQWqkVKaEJD26JM4MDQKArzs7L2YCrczqMpuNfQu8HK
jvkjJHMi1dKf5OYyyDD5stmJtQMJjFfUZJI8H9kbuJtvQxqg/IXeP2qM4rdyqCjd
wZ0KAfO+DgWD5qJkj3Z96q8Pl9f9OBq5jQfQP0xrYgL58tvmTnP5iX21FnpLcRnt
nIQpj0acZkCz4RObCBjySoDhg6KCXgtg4PRJJ3vpw6PHLop4rfVKvpbaLJBbBmwS
Cbu1SWnPu2GTvB/CRvutxtEZTiMEXEtRAAdSnmEftAKnsqt3YXHKNrEJHX+PKjHl
zbuj9q1ZpO1d+kKjPbc3C1gqbAtGWQ+r5iKwCa8OWXy9FIQQB73c/YeHw+/wXfCA
z+HKvMGmIKB7cypwZQx+zbVjZbb8Cg+fZoXqBABARyIdwXcxrirm6NmMLggC17Yp
J6liH72abfqFGTDpl47Wm16YVQZnkkXgd2nJPf3qklZsEQT9Dzmcjzict0wH9R8h
NreQA78ttdoVTXAhCGASnrZwfoiwPtk7yC0kv8ZW5ShUffd1cH6tpb0G73mZa516
P436boMeICwgmxs6Zz8AjjLdt4pAWNjv7OVEJTFQXodOC2l8nG5IHln/1vwQ9lNU
tOt+mGObBOVxwSb8gM3ZZzgK1vw0u8+pWQW5MVYmfJhV618jTklVSkFBUu+NrAwm
5byl7N4OyiIzRpqPAuNb7zsMU1VoFDnd3YWDaafijfZ+O8kVFjzF/parwi7Qydn4
8Ek2JkFQRZbFoO/ic/4UmxJKT6FHZ63Doh5D4UNqlB9Taxi+EQXeh7pLaxJ+FqbF
HVkBgG27AiQkxfQ1ySMlJ0MFvDDbPQ80pl5OWFFieIB0ukMzwEVf/4aWc51YFWHb
En6ELLbp68+0cNqR0DJ0ckzZZBkGDSka2nrnGjgiSPqryLxmVXT0rs3ZXst7qGp/
IbGsi5cLQWj+93xCI286Hm/yko8A6xOPwSnGK8t+B4qqNNpxvLDtbQ8uADa4EmoH
sRh8yNE6E/RJiqXUNLJjrzpa96ih+oXxkGvgKllDFP/lfR4kTxgb4m5IsX64n+9h
y6yrM1DAh7ceYg0/SBZvLr54ye2vpDl8TPEF37CYkpC9t/04fYS2OdcEnqqmuBWx
/oihl/jEtg+UZ8t2hVlZAiz5C/d8m0fIS1qyt6nEalgDPimbkVVNkyaWsVQQoD3Z
p5SRHkhjLkbKr0U2dX9NznUfZNOCwlruacyAsFsDM4XGGHviTAp+IMhzRvmSF8md
M1sE6BMZjDgQa41quh8rJXpWJF3QzXW0EtSEKYwdwemmPHBH198cwYZkvjFuMgKN
IWMzf8x+EiEZxpXWZgtw3PZuXGqpjEpJz/OJ6FR0i4oZkNL3REIdhlBMQMepTPsG
RxkGq/vp2gSdsFNuMidm1hDLiezio/oYgnaV45S3UOYCaZg+JvRNqG3ekVIVbBYc
dSmwVC6NnEIXu2s+nzihIxkNEkCj/RNqK2DvgrzRR5SrkOYThhUSj1Q09xyItoGW
rN4DLN/DMb0pm5gvh8pkM4DkodxuVb9MD8y5j0/oFXYJkM1s52PUOUPsN+wihs40
+p0WRu3uvRDCFqrsdaAKYFrGhF2pPEvzCrNJ9SUhrch4XK+p4wue2nrGlbJBZq7N
m4gcqVMDeOqAm+F50yDjhOUyMOKTipS3Z7BUhN/MtVFin/emKHk5thgnrnXrQH1e
P89UVCvTOT7NvTxuaW6OszD3grTj8a0f4HvTdEuCAk4Kz/xHP3gcaF2UPSbVyPhG
0MaHitxltglg2YYcbJ2sTBn+hHUEhEsdR1gN+rVn6dXz4w6K1q3g6YEUmgSRamuc
zYycrPbK3XQI+Mq6HJePanp10IaOqJ1WdpMIy5/p9yMxw6YUjdhba3k37Iln3SSL
sa0Y4BYMk3lk5sIN9ZxUY0mf25iTyQUvhCkF1GfQs8M1AMajWpz3kFE+HxLJmEUP
ECzFyVQe1titcKL7tsNvUQhwfSgTzRkdSmulEblNY/4VBOjwa7WvxiJZN7Hat5el
iI4j4u4UmlVdXxRM1GqF4/bvti0C4ixmxOL+n65Of971KOnGCRF/hceBNwT/G6z7
mStE6fOD0M7ddVfvtPOEC90yxXeiFh+VaFIx7YBriTxwb2nNJSoskiEQvezJZsKo
lpH+Car+o79HAKMDQcEHno/Gry96SEm4apWmtV0MQQTPNoTqX3M9DmvsaDQl0Qf8
cctoAzKA3DX8MCKZwblUb2JZ3P98seaRByBh90U+MwZIFVDMrVc1Jkt5y7q9jBuB
Mdtm4K3Z5ksRwBXCn1kx2N+fsDd6UpetOjwG+MjmzckkbEX/eqlhYPU53WtlUscE
fTxDdpSkC0qELfr2OWioyQ2g7NoXrBV6mvyAlJWFkfPZtxZEICil6v2c4QJi58fB
8VywRIDNvEzO6NPTRcFQSFW1pbC5AIQigyIye7JBTCvYH7cbCLdtUGrYn2hNVzRC
C+8hQoptHedrRdDhAXnI93aLnRNkeGl5W18n9+BKT8ztplC1fqNeHedaHwImlY37
jvnpxRh3UuE/4jX1pWaLSIEpLOn870TjwigNQ1+F8bbrDqkFCndfA3PKKy+GFN6l
OIbf/tSxjKoKNyOnPicqiC0vGrVbhJOBNGmrnWZvaulTOtdSfBLKsSlBqPf/Fsfe
yK9IH2ndA+IXXHV8aIxoXsJG2Smv5O3V5OHq1C3Ktz9YLj+txiqhjjYYtnxEKCeb
E4i5rh3ifQ5Bjo+dnr/mUnW87i7RIuH+C0BhfnnhO3VhYyURvLFMas3wPTHeFBxj
KtgkaPrw/Cw2K5lKsYhQcPv85HzPH798qECCVsOfVnA2f/Mm6Wo6DrxhCQ6LT9dM
s9rVfl++vFQzWGPBN0Zf81TAGk+3n6Kk6uzBaLxIcYc0OaTzgfFg1KKToxgaqgqk
TFkP6dsVv11CQ4XP/I1ehMTQ5E7bgOQr/zCJlsja66rZgb3qzkJv9aEDLC4XwDNj
UuJx2WSGVm0TCT7ivk2NrdK9joeZmiEyMDOQfZTPgfJnSxv1CdeGnAaIHMzxGIUm
N0oej7xeex9gWaBX8iI8j2qnT7q8BqYJPvRSgQ4KlvrducZacZ+Dyu5jW7AQMld8
geVGNAclxSHxGBT9PQ2dqyzCnmO0VGg2zVtejwHVh+U60Rl1IxD5SiN6x0c/qxDS
4tt+Oop62AeGAQDk4DzmNN7y0MEk1ZYuKSrZPKsN8rcJs8S1pNnlrkyUNdAm3P58
6bBDumcvb3KWDG8Tx2o+ANLyq3A07wiwwnEj9xeokGSbCbjIr+OfxPtG2eF9+RRA
rHt2+L61i8ZU0IkiGDzs4jb1wcu4sN5c2MxcJbkgo1mkBLVBjbjFQImeZ0iSOSzF
kY7Bf3KENChA4ti4/LFuNhVHy3lihGIo7J3fA9JlI1aEUNTnwiOh5nhAoNdUHrJh
2kdTQE/uw2dZC/5/Yw2H1WSK4JcxRoIZYmxEPIcfV6QARI5tIu9NkDB3r0av9xCT
VZy1bSFXYYqv0QDv8Nhd2WIkCxsLd1cQtQFP5bOeb/ZWDD9+oUXoNI97HnJ4NK5O
FR983ByMsXJ5//wOU0uRHlj4kShJTTXCOd3R3sDz0HCbhZJeQ8WUQU+IdqfC/JjH
0008MGt4vEdwp3Gik65dxRvMdnXEUvsyz47H3tl0csR9xcdGyZPTiI3Y+X0E7Wcd
E9m/CJrDS/INziyYenKEegMXCe+DogWF9dnjE8CtvAQ7W05W2zp5MTqxvgiZKEL0
rCTjF4qtGZdESDHkPOLm9IfwDnUHSpEAVb4YCqWS1HFaOFdJFaNThEsLbO9xDqYM
/gNeLO5E0MugbBppVvvPBf4L8ngDLGpyTTluWkrtyoFt6kkpORfm9jhuyXTP7pa+
aDz6GqKzvUtfYNfS0Fho2bD+R3VbKy80cvfjqwjz+k3DX1h7p9LGqeyVjFeJHNsj
R4BjOIJhCxKaHAKaTdL9+dLg2rFPaoBfRHSeZcydWnSCwQVkYpcrTIE1OH/pr/Hm
4HXuHDKlUu2EWiE3pl5v2Z6bNVeAzOX3Xnkw+UO1AAQPKx2Va70lFz7b4RFjc9LX
hdaohnxl2Xxv/RKHJq4IvYU1kL/XPJZ8dmy6QgSnaLvu+DXcdkS6Kdlx4hecqsQJ
Rf3ebD/XrBMIMNoFU32qhlYmH4wrmAP1COGDWf780PQpQ+s3QmYfuUyDMO0VWFAQ
NF4XnRu97Ht0GUS7JH5sD7bTX8ABBFR/Cs9UjDL6FGOmawKR+MazRjPwnq/kCzIO
7g1xC2fDRxahBC07/uuSRwpKw1Yud0BOT4EO39T6EbUK9k/lLi6qIR6SalC9/+l3
SPFaqkDnm1g4T1bxdvbXIkTc40ha4Gq4vq+hlB8V08y3OEZbFp0leeZ8NEhLUGIC
hmVadpcwOgF/JCiGT+01p6/8t2LSG0+xcHmHlngiCnh6QCaW64Jo2F6sGC6R0Byk
wOhLJq8C5Gi/gR9GGUKPOKBBy/6ZTk5tT1teFjBNy7tSDyl/nzPxymZW7uz5DLRd
SunMtke3gm5+2omNvnZBxWpZoFhScAOq4QrD+UYypfQI6H+GmsK+7zgI7OwX+hgX
kpY2q6oTLHw4d/MwrjanNXxjAhztZY4J5vw/0rhqkaLPpTmPJOdjdrI2dhIuCRVQ
JTFIuFVC4YZL9EWKf5y6Jv6AYCRWEAjrZiSgCLrLOnht7sKPhvI1YL4rEOlninyx
DxDWEszn8xMmyr9oIKlC0kcuRiBFK7tH17roELUADq8mty1X2Pa9L/BzLeYMQ3KM
cK6ZYVQBq30dGGf4Y2HyfPAhV6+bC9voH4CjDH151qJEew8tM2ltfIyJLxnrO8lu
vPXjVYML0J++eMvQsoUv0+FWPmJ4jmNyDd+wiuFrKNN+huxwxRE2Swq5RZXXMcEs
yU7haRel0UhCk7wY41V0vvhJo+uYJqDscc/vMHWgpMOeAph7UzAJ2Uo7NEG9GJSf
CoAAgBc3KcMI/v/6FFaB8MUKf7hIqSTVgcFmVgkMJpwIYqQL+gO8Qso0EFO6tiS+
2L1DjNjSA6EYYrQMFeR18YAbz05o+yu688LZoKc/LdxQyeClj9cyE7Pp6U52KuIe
zMeLIZRg274ES4tXlUe52PJ+KDFJj3eMzDRh38OtiueePz6SsoabtmfvYqjd8pJU
6zZisLgKPKiykMQsigu7TUMsVtoLm2Q/MDJYeL/A28jO5TY3oXOETh0echlK5fgN
iptdtpWHWiCkvky0PCtAch3vZmjoc+8HMplwDven2mjaFuEWyPQFI/eo+rbxetDi
QcZpM+CuIFL3x6igkTVJQRwS+FkACPQie/XHoTSUYXmFQ19lI7DI2Nsn32bvQ1Nj
YKIWh0V9ZH1Uuv1DMHIeFBSlfsmJ+JYGrnoPd/4bJVM1yzAqBe3deTNB4lSVPPEa
ashlWt76Fe/rUKmqv9y+9OUfWWl4YK9fnYDO7XDzqdrkTWRdJz1rKpo8KcXo4ntP
QyrwyGj0M4SvqxZv5mzm4umbLJQexLCjds0Iq90Dp9T9MFplVL6PjT1Ix3fV+rxE
cVZJBhPGdADgDgvRwAL7YDVvoXnRArLQs7Zpm7XiJ3e3xGXyKxh1iuhpEJdvqjrJ
3kTlBoJAfQps5/RYs41/7/CiQuoaF8mocULOKx+Usc01tJX9uTxueyJP6+wGOLD4
ZnZBD40/XS8tWx5C6kZSQKZmUhCiDDJieUrPQuV3OucbOUW3aL+vv0u5u5XARhGk
0C+m4u6w2A3L6nNjMnQcDHRAC89f25kv1OkyV4qFOxemEbwLCTF7TD+FXnJJBcZX
XQD6ZetFDd3j3POYZBhRY7MGzv3I1M0uaMqHepv3fFGP0nJfGc5TR7ZapzUrAOf+
ZBlEFCZLXBXTjlOLnKMtYsDklYzKy0QmcZUC78R8sAdzdtR50qVXQkHYy5tfzIK9
hsugdiPodF2603EWryhy2tf8+tamUGobHuP/8G/L09UtmpqONtpIqsKO22Y66oAg
x62XLwrQLEKqOS4Q6MD+yRk4DYlC33JfVBqlYVekblhC/p3XP70lWHb2nnoJX3Ok
4oyfPEAi5GNOoTZxqOjtYW/w9RgH+2/cy2IbkwuC2OWslWY3G/f++8iMwdDCu5iF
+09j67lYjYvHF/0wuig4+nmkqUYI7DV2RO+jZUervi6NHYgvMfTvXp1GbC26OtbE
Srircr/YDrsdGqW5MywEpIFLnP3qScf2ln3MueJpj//Tq/Xs8ssNF3l0QrrnVuXh
gebGB+wXrfl3afyPCFx2kCRThFnjusurV86M8Iu5Ip9loPXgsLXxtvRuL/aWKgjM
mkYRYfqYkv0iG4KPPpjr+Jkmy09aU1ota5zuit2AwTDQoVld2YytkZW6EtKaQ8iw
Pc46GTJySXAl+682sPW7Mk3BPbf2CnzA6staxRYrPdkL7d81/l2hjKEO7dHQz8rM
+gacIWInhJf3TzFjjF8Z1s/d1AbYzhbPnrdj8lyCoBY2Cfd2wJAtO/LRJtLfX40x
IfQK4GAI/AHjftpG20o77mTbYbXwT59rr0qc8GHtam1QO+qWFMSp0NnfRjRlsE5e
AIGxkBBsH41Bh6ngtTd0okbJgJjr1jyOG+rgwEs8NC0E/Pa2JWhvBm1QckHpj1PW
1F5V2tZkddGw8PnK7SXaUKk2ifQGFkDbqSDcH91MB4Hivz44Y4NRgretP13dEO4N
oqQA3o+vrAIqwwMV04tE3oCQB2Fz2qJTWqqMxLZpo9MU6qQkv0G+XqkWb7FM4hlm
+3Xbsow2/5JfEYjGTBfREPoYh25Vm+tjY9hI0fomVn3KXoa0ByqUqmR6sJz/P9hk
v4sXitgklhpHd48NZ/e1OFDygWiYSjFb3jUKvWP5Dg8sR+CAfD6FpB9h9ockJyWX
SZU1tQ9tnaA97u2w2ttod5l6XaYX5sNEgmJvO1R3MG3H9gElrJRmQ4HWs1r3NF/Z
jr16wtpXfEn/5H6EhLOhaHPHK2PR36gXV7Oi3W8PfombMrmjxi0j1kP3Ne3juEYL
Gfo3STJpjyNrKPlaVwLrn+2oKLXBEYLN9ULkkmx1QUs0eSF7oUN5RTzXdok+9EcI
mULgyQE85P5yKhKxASjJUT7b3BS+qsG+74kS/vJ7rbeTpfddErg4l8RK0NPzGMQY
K2DON3rw5pygltsy9Bm6nhKCOEVCmR02y8jidTmsjcX/lm6ahkYdh+qOFfELu+Hy
SQhnM8WGl6rJ8K7hkcYwJNFLNz0W4latcqAwpP5WsJBFbRmT76uMk2VUHAo6LHzW
YwpDYY44lGaXyFMLhV6MI00mnh82RY5zxOsGa5PoJ9kbP3bEXZORkgSSAJiTGulQ
DZVY5944AbZd7RhHqPg7/RGIeIHLxh+9LXr3xzwZjVf1cU4Ss31IRimnnTW3RQOR
LRGxTa6P2SCaHBoqiBV1fx8ABb2iHxXNuIZ1qe2MRTiDc9Ldk3EiH+XO6Y2Jue2s
5sOp/vwKwBk5gJkuoRfqW4v0UqSl6afg7tYF4I2m8cQf3WpxKbZMO2etfHlElGIn
gNoS9lP8zyvBZN02IlCjmB3411N/ed/aoKJO8WdVNxNOrJoBilVz/0/+Bjg7kdPd
9Pu6qK6VFZZoJc2V3Q9TL9qS7Oj/kQzPDbYYwUufIv00xuMpoQwQIrVHJhdhs56d
7+lMPxLUL9ctmPbbjvAfrqTMzAwWHGIVjhHp79hfA5MbkqBLrk6y7xwUh3JmesXW
e3HDfJIrTEqh7BjMzDVeOGjhncKMR2LX+3ZMKJ8xiSy4gaJ33ScJWV074iwVV6dp
/eOiTNv79CXNFmO2zkFg67FT0ch8SNkQPtvXK0Kz/LXk3zPdyLDWZB8T3u8wgIzd
SZfTwjy78l2wLf9BKr/2qcG8rrVMOBxzB+LHYY3EUZgYfwMdCkARECBM1Iz9B3TG
w/wg0z7xahvr2BJ8px18qAAk+WcSnuRbeDN9xQx5zstXlxPmzdxiZDg809zcXr0b
m9fuRiuGqioWXMTbHLvRlKH7ByV6JPoay5gau60qTEiq41H0k25CMHFJF/1Qxo5t
FJd27JtdS165P0oNttk6B4qXW20YYDB57OYQwlYTB2DBTlaPi9uOMWtaO0enTnW2
LyT2HeneYcpHOGKnM0aW9t4UU+97masCqxm60HoAHei95URUEqPpP64QiBDw4btf
9Iuo2Xfx6TwLBWbUD0ngOHz3DAZZeVXaHtq/lSXP/U2MxyL8isJOgF6tEivgCG2x
uByUwzFPYahisiEgq5Pbm4ueFr6QkuEwGMu0tKZXBY88mVX3AZKJoh5/YHinr4Jk
+4hZu9DqJYIofJnltPt9n9E6FQjqpyx/QfMzShe6TIlfkyQBn5R06AYYcSLzwFIA
NlO7PStMUdi3gO3RUlsZhn1WURayFqbuGLLdkc09bI9Fx/IHSC+W3ugLGM3eZkGS
1hlunOhjKA3lYatiWCATxSFDg0E/x3m6pKEwse5tQTgqem6rLGTKb3h5AgJfr386
lGJLZS3Bm1CQ64TNfvr9PPfhKbjdZB9MXCRjSTsSllQL4HaTYmA9xJ/mBrxXRKl7
ssSkNPH/F/m1VKz+PWvI9xouUxlPPaPoIi4aHqiUdkh5yexEbCaOtbWJ00WFm+3w
FIwVSkws8n875+nUGP2X+8PIxwuiRXW1XW1RYqPZkmOC5MhGtB5BBW2oLHdzuXjR
zYLiJFhRY264PglERhdv/uvR0cQ7myE92DWhNj8Lo7JmM8tagui0htFQaHIYY78P
YFZka93DCv++wKlE+0LieTZxFmhDfLy3Wp3+D57oU2xEhH5sEFqmWEs1fLSHiBcG
LjvrK/sOnDMp63jTd/ngesXEp/MaVhbq5mifjw7bks0UUeVZzTbZwuovoACxoyGn
mLdTo1cXixUFkpHh6SkydBmXe65Izsue/6fm93qReJDP83OIWFGuUHSYkRMFv4QX
P7AOkxh/fUTigm7YyWqEJ5dCaIA6ela51BE0SrG9ebJVf+KCjsh2X5OhD1mtKGtQ
z4cNqZIWsDWNyjhrm1o358szevm8v9vJkL2kY4ap9R9jBTafWklTpped7JyUpUgK
MGrQIs5/FyghaR4gzla8nIDGIedCMyrAY6oxvNoWLvM77WsM6K/Cv2adwAhirQHv
XGbjlGXQnjV17Z/mlQlhwTcUkL+cHkNEaQUXs5AjZE60LbzQkD11YoDjOZQDzlAi
QJ6q6mwOPyPdW9gX4qaTKa4KFiB4nICKoXYZclvxDkN3AZe+sq9cRSebhmZdGQO8
36ypm9z9hnEYfRZUFElKuVSrrvN7AP7dSXpjBlsdV8swqNsn/mnaHzruDQzUKpA7
AKPsEHM+kcUbRZ+5O2RCTtT19l/KafmT+NK0IWLSd0iLFSnVr1+FpnbHfYzQLnGe
Ok1rReAwuTGOfZxJ1lDvWDg2PlQGHcUz0sGOMAZGJJjMM4UCjgYDJQS0/MUNjrDr
Ls7BGzo8O1bs2MQ/M/9gKBRyy9PZdI9O1nScnlwX56zng/3je35zn/EU6ykGCiz7
//ZTXLg2o/l8F/OGhV8DgdoLIrH2VNxz6dU7VgaRvF6LgGlCU59cPz9UzdxxBiVM
ZsmnRM75QPLa99NvYz8NfsfQq2LZUk4p9++Yju7Qce+npVRLGkEhNH8Rf80qCMHv
FQtkfSM0QIY3fuziER6kFKL8SARRh7fD2HHli2pZA0SUKpyG8zXr7AZGK/Qy7XP1
ica9TpBGo6m7BVp0mXlm0jt//scGBAhug1W3aCTKewCanAPTUsQHZUg77ORYXm4f
V8T7kgCD1RhzUipQpnnksargjLgyJDemr5rhFo+mRFJLxaEhbCsfMiwm+qWl7A2m
d2US5GIDkheLfBwkkhhpmVVZ8JLcXYp75pibdD3mal75dSLrV9oAK/ErekKCMKvL
vAiJuYZVAqHdMb+TgiZbvzXWPE7BBAX1jGBR4wkHoDI+6LMVIVqBrfAuWRkuQIUg
yT+rzwWqyj65K7+/BhdbkooDSnwWEfBULMxJ4FGoqAMIDG+ecxPhNoSGP8+bFvpq
Y/YZudHoFgTEI/ismaUXOLqnIQhWjoODzTS1n8xRAof7HY3MhksuvKp7R2lZgpOO
IBK+6scvjeeo2FVGHOOkjPHkqfcVy6nrEPBdtCtf/mfv5I1WVb1vX+EcPe2a1cLh
hwAoO5DNFdvq7PykO1JpIyc3XesQAt5o7jlPYGj+1gz6GB99BW5Muahd/sShVz3L
qNtVwYorVFKiSTfKzKXvLzAEoOnegqeBQotNRM2TqATrvf41atxezF/5lDBNtxCM
GOcxYkaKGsE6LsMAZrq/Qs/NUbt6J0fbfQF0oZCIM/PbocKvy9FtqRnasdOr+mSf
VISr38Z8ajhCfMcSw6xPc/67z89llzIN+xUKmnpzZ5qO1H9sOLU1awNPcaGnpl/1
Z3YudOW/UiYaLP/FZs+56Ju/Fp+IInD/jFutgEiQHrlEu4T8QrHOgHXsfrXhflMN
Sz7vwujF/UFf3UoYxl8xBUc+1avgFAmrxnMnSTaPXBd0TGtHJ1XOkjU0+tjHUPOr
DGqM9Og4dy6Iky4yrQ5auSm3quQx1b9XYeKgFiVH45Umoue16mMH5tijO0RPD+W6
T3peQ4UtFMff54BR45lbPwzf20/fe+KFEe54skUcCU5SSbWkTByLeww9MtVPmm1J
jqnjRtTb86+CfXISm6m8Tcn9CYTm6Kl78eoyFkFD7Q9SazFjjinkmFDg+4AcbTza
Oe1zkaC8Kg0ZTgfr7ouer8cTbRDq0xt9BwMV6v5gZZcUHJXLuBNUhKkWeNekHd5h
UedtFWb9cUQ27DfBx3qtlyIuRFi1RJO0DJ6qY6f7iKy6Y/6VSl7pCKCI+5jgzkNy
VucEAwffIAICbCZWA7EXi4urdALL9D6SvT+kwYKNshGSw+LP/wUnTO5Efs40rHDn
KcLj5FTWOhiyT1cNPL9kgLMa28vpmoi29rz7KPW0t2PU0vigPQG8/nI2vECkSyST
YIScwpmAZ08M1Hc3dOtKH0Fd+iqqtao9abuTOLaQ8m52B8y3SU7O/8rx68rSGV+B
iLNA668610EQQWg6kJXIiupt1jEGCDeA2t+tFGXO/3cKcA12yYtlxQpKyV+ILcgw
2RfFq96EeLqDp+8Los2/W7vkCB8q+gOjCduDgxIpVbZlFbwQeBqiyn+yTufwMxvC
gh7VOLuVNcSMotAfR7ytQn6sgTSrGdP4ulgmKIyw3cVFZuH2ckDqCKWzkikoU2TJ
RMwjyrkQnqAyL6FfK13Xbh3lCyc0jX3rm/rR9FE1zqS1CLo9BnJMrDq8fo6zjOsN
y5e8etV/RPybrUGL2Drt33eFPwiO3XW3agKjoT9xSF7CAU75EgzzJusWVTEUUkWs
nTaBqezehrIB0jPmDLPy8cf9cOui5zuxF/i5q8AyziegMwZdbq9v7uJkMsUwwJV+
XxKLz1zBLnkv45g01S3KNZVAulu92cWosem7Cq1ejFQDNU2R2T3X/cc3G3w41ZQB
sVpCauRhSSCzI/n4MlSW1tH3h+qfrh+VZlDw50A5+EMqWw90vY3LulcSukzIyaf3
cz222/MNdgMoimotCYfRw18Ld/UbGlzfb/usAx5K7QvKnGDgLwexMIcgeALQv+1Q
QxnpkQ7C2ibJkCdpD9XBAzm5K8DatTzSPCYzItubzY61ioCfsl54C25xKM44rUxt
JgTiLO+XsGHzusryCTw+wpQHNwoWnwVi5AvoEitkU9n9YLso/1V8Gp3DwCQ00bRj
V7jk+xz/IBFZLCSu7alH8BZOEfIcm7jfPj7693yXuQP/CowdY7cJhCX5FxQDoz5O
v8iu4VM2+klC4UjXzZwkI34msdUWYGoDXhBurDLNMoPTCIE/ssUi2PTlpR4eQAuC
JXYQpLLLPUmJW3/ixnATCFV7Fr+10DsplKI/tSS/m1o6HYvtCHZtGPKgELtC8IMi
McHC60ZsMEFpsPEvgcAqu677OYDWj3agy8mWNeIVLEHE4b5KdiLFQbz8kZnK4LEe
FzZBSLK/b4j9hJZlksotEbWrJLVr80ZNd80IWoUoDgCMIu3uJD4izUlK0xLNteY4
f/BVKxWOtXneqkEzf01Tn5jZpfaW+SuxlocoiTXGmr57vbunhPmNDLNguKXHHWJF
fb+tdcVMKN3J11uZ3zaML2H+0aRsfUM82yr/IEyIJKOK+kLZU0z74+iTif5Fgu4Y
D7rkobWJmEUkValcVkWnC+e7fMPoKHdpn/20h7yUltT1PZlNW80yJ2EPWwBVpUcG
tddcPgOl1qQjR/yXAHPcVPEdYbMtrqgeOZaBK3nLEZnCAgvbUK/rmL7hipd9scH/
BOPXaej8KTjaNpmd5ZQ/Cyb3UfFQ97YQMoyb8Ewoh39CqT+fzfOnDXtJBlDlFpZp
LUEO5Ij1Mzqq/CPgm6eKXxmv7sRAh2UsRXg6jg3hwmF5/fwaDFbuz8Fgpsb66eq2
TZItdXVHNvO53Liw4cHVmyeFIQmEiLmPBM+P4I1O/OVgJUPdw0yjcDaxRIv57Iyk
7J3VRlu1LAEeHzY6MzPvApH3zGxB5DsjeR5ttoTW6QKQmGTXm4rtjZov2DCfCwop
CZGuEbRJGkgLup+/RSlgcY/Au0+sOsqpVvNHip4O1oi3yMbgzi0GFkwz/7MNRKeS
2trTfQ2+vJUxwHQiAw8kvNYWdlPYGQvwL7qn5x5N0rusyDL9Mx9Dp0qDyoyM/MGb
u9MY7wK37IQnAOjJeRh/yCC9sIq7x1HGwwqjwceJCObToNWckqB1x10+P40gjHii
wx185fxTt/U/ifVlLT3G4h1gqsQbp6AAF6eopqwftegiBxdKXNANeV6/06d5aBz2
CYuYCCJrHCMtB6sVnzXsjluVQwacrFQxrSuvYmTnURU9t7WvMIERntGAQJ8c+RNJ
rFN4c/ci/R311T4Z3zjNCKjHcVtP/oF84jTb31f4PX2gyC9gtPe4AXDPF3/039M6
MWPt01bB30QSHvWHwsHT73tynuttCI+JSPoxz+F/0pJt1bmTQxfKMkIg8ciaxN0Z
MJb2u7JY7uQX3ZhI5Xj4vPlmoyPJ9JbXrHSTE4UGRbmfihPUIhJbnetIYDZQnJYf
8QNJs8mfjNo/xVy97y3Vn0n3kXPgd3ELAH8GEXQMiEZxUBuRp/6BCs45eyuHZd1C
pUZA9GORxnAZ6yqHic9HafQ3P3u7h589yqkX7Ez9o/7vzRzoqGtp2Nx8KR9wYMfH
5ZoUeEwDcpTvcGl0VXzOR0DGSP8wsgor3s4Itrb+9fNqmbvCJ3D8M9jYFKORsykX
Q9i5usPXbha2Um5d6rAVGGbHroGM33zhartXOoK6Qz47P8Eq/yf3jER5rEQO44xM
IVakEQ++v7/Cc+VkWPfIF3xrYIIzB9Q1cqilArBmT5DNFpFOrd/CGD9vJCOycAak
e7ZyPR5CTPoiEuX+pAr7/xj0flBy9WsKpwXos310muE/17Fi94k0Ffg/xYGsOodI
O1grf6GuAxjs8Y6SbgzT2MHgcJ0xu9En3HuXuA5r+YnFZizYiORsoBe4rFGnaEa8
rxRn9CVRBdgewZe/EEP7oSFOOYLQkmW79TsBjYL0oFvA3lQ59Hrzn7xfYpDyj0RZ
rSe1KFqsh1H6rgJpnsQQi1cvua4/AqQ2RbwCT7/hrUYHRYQYpmdTLURKFzwO9h0I
E88gtG/GBq7q2XzOpAvKanl30Vd3ac0uP+QQjUOloz5Lyrx2xSUM+ZPfIzeaCnk6
h/3c/n8MndDnOjk6jooDM5HcyDYHQk/u0g8Gp0mQmkXjNs20DsrBFhIurkU4cxzq
2wUu8QB8PNKPpb1lWoAyzvjhaIvkvkqOSGxxSTfI6Glu8nbXH1ygvYTnyy/rL+fC
pc4+rC5DoXiIi0psR29qYiNHQOGNBY2UeoRGUqcNOPfsKUicvf1Q5cVhsaC8XeGd
RvirrXwR9WNZaXI+IrKr63dA8i8pyxiqllIV45EU1adzmmfKxpUJYEPcPZqNYMYA
KJ5KrU7ojnN8/JtTbLDzRRkv5Yn58jTKsEUAqWDW7NTOBaTa5AXzKxY8bEJeaGJx
VJSe4Auy1RFYzxQanHpQVqSgU1tbr5H419RgMKmjYVYk06uZvP/jXswDN5wvgauZ
byck4Q4ovlN5/HleYUntyrx6eUA1oyPKPOztTHD2D08Y8IMTs5fxdOvf7rCgPf1/
L/IEIeu4R/npRCpu7qsiHYlW6DI0fhkMqF7Otu+JkFlZcRDS2V+v9DGLsSb/L4Av
pS5YEG/m4a4dNPmDW3AZgfLRvintCY7k9Q5UOlfgTNMd9fGMIX8XQkJfAwdwzuJx
koAkCgBEwaFMBkGtaEwxiT+i0Ek7awSt8LLSTTgp1mO1McURrOjIBVY32VFOZZa0
p+F1UMsEfrTBMD1q1VZdd7GxSI7/PQF1OTYz+9xa1H64LYHJqz7+I0ZTSxj0LYcv
X/A5rzsr3BSGD9TQcqDvMRMgeWxW+R+tyQEy0MK9Zcgq9+PVaxieLSxFJxAO9rac
fgGEQgNB1KAuhOHmJMq+ykzsWYFzhBIkemoPR5WehT6wqFsOI17P7avDBSYy8cuS
sxPE54tPUgBX5167QWSFvDG7Cjz0tTG000InKk7QLfX/nlPMVoUZHsfnmn+GYbqO
MltmAlL1T2Vrrgss3FhvlYCEKbP4+L6qXi3cu5RSu7fVdjTMdAPdKviiuL8WM8Hl
7xR4ZCPlX/06Wdwtgen/FLROMcdnIlSDSTMzI4DzE6gL9ryTmKD89IZfMjy/+m4m
ABLloVruZnFaB9/jTUSMs4PEWDQLNbXDhjzgXrkhUgPfX+4G8l9jlnEjYqilfsW+
3F1VxX1mVdlKWoWtSasa3Gt+LECO9sJCxV8rrkpeAkfkvbtTikrYcLBrbzsHqsWi
bKFLukLH96XI/wpd03PRtzBPtxvHCbePl+Z4XOWaGnlcN/cfrjKjzvOTn6SMPQLU
650yEqpkZiqFlw5XhGpKaCwRNbT1TKmvU1X/wRwNqWsRei8TVKpOpETqOcsJVKb6
rmCbxVBHZx7KL8kOLC0k9EFrpx9SvPkt92MIhIQTJSUvoWyA9+qVtq8j7x6ap7d6
mi2fYy57AGK9u+bmFQcAwZBFDyGmuSSRyG2GfAxBGwO2E4KAlfn+RT8iacsqmdzM
xxU274ITpolAX6MGIiohpo77BiLKTpYZ4CAFCtuUCt7qr2KEH9Aecx3zjvCdVp7F
PL1hXk9GkM7dVSsRiXnhQ2qseKLmLbPsTxYRet9+Y8uSXBDlLwxgce50siaHSDah
Xz2GrmbQUruZ+o/yNs7MtHheqMBV4NKF/7IlDSAKlJ59C27NWOo7yJd1LxUfviVB
Io5j7DkixjGLDODt2NTnpxFSc0rYo4UQ6+7r37bNNWBGZIktOGjnKWiORZfqLS9Y
Xu5WIXW3mvqE79A4AwG54OAcqSwlE9PFYLgvZc7w4ApVsJ4CvY6RODAsjYw371lk
1vkCt31x5YjIEVCvPLYFiMVQQt2QzUhS2lStJrdKzUd+Vh8g/8odSRl5ldSCbJ6l
wgMWbC8k3hL+mn9k0A7uUZj9G7uHxunmC5Imfjq9UF0GiG6ee+H9O4gz+5LXtgqb
1ia5U0KCEWMHU7lCSAJsJyOo4GHbP6q1l/fYvZ+skHF7+mVw+dI+BZKGYbI1RFzK
N6/F+7W1weEWmXb5LBkwctlTGF+Rcl9o+QpFlC4sEkJ6vFa40i4dcuN1puax7N4J
9yg50T3KAKZYqIfsffYY/dvgPYZ797eLPpEBuxJxKrb3BEH/7sa4YhLUMmQYpeMv
TDtBiQ8L5Ibj2SSBj1fb4lL1UAjauSIuG2cFXiuFs1Q0iv7ssyYr5/Blhrjr7DYL
b864pUKd+du+lQTjGxFGNHFdWhrWt9lutfebywntg5rcA/GQ/GzrFA873bpaBGXG
3Gqb8Cqt2VjIYYcBn67mt5sm5BenMNZniCPsZdeTDceU8g7OBri252LqVB2IY6mE
IQdj2XuEVBCJgDh3xpGRVkrca1GJVytb9DrjFjsymJmW18Xdd2kmi/ykDrVAed78
0+rGrS6he8LGL4eThhUsI5Jw/mAuna0VUINGaqq5GxfDrMzcbQ/iqh72VSpz+Tjb
PbP6m8T1dQrQ/69ig16vb1Gcm+I4sLU4e5zsdsvr1dV8Cik4zf/coxvyzjeggdwQ
Pc2kCaneb/SO/dUJ2y84E47fk1tXrSISdQFdtQVVP4GB/ch/Y0OaSeS4xKJlvih0
hKzSqMLxIpGaUFcQysNrmxzru7puKYS2PRhM3YzZfjhwGus6CdFFdnU1M9zSQky4
GOwkNCbeP7JNiFHOBughEtDLB1GhQlgg9Hhg9Qte3AzS9alyuh0iYJscPkJPerhx
zF4BKalArh+53PjOw3kC+G7+NHUWgDh44p4FErsPPY8xc7K7yHvYEy283ByZMDPY
RcLWebpVmNxrfA7wNisg51xq7SM06uU/FWXAZxG8r1D7/tCMOIKRMyk2/AGl49V8
091KXFYdhKb3FoAf8OxHOLgKVY0iToQ23zFBHA+kYQfPorjSfC3hXHW8WLWKpJcW
Pbu+P4+8v0ZTBeIpyVCkqUmg6EZB2gqaXMK26qE9o+GYKFzwUnQWHyEmcPMV8oay
SeiFOWMjspGuo6O1HJuWYK1Vx57vkL4TOI1kc3jpEwnGwZbi20yppv9nP4YeVIuc
EO2hE+1w+DZx7kXCGSafFC2ETpKlaz7qerIH98cuLCcHaRdZDIhe6xyX0x5LOPzC
5Ip8PBh5dLlHepHwdUSSlwdk8ILL7ayieHRqCNFx8v64t0fOqxsi6Zk4maiiUBck
Z4pdguRcNO5UEqwAJ1LKfClOFw9FHvMHcBh7Zv/Lp/zy7WZSDW3QBUEvOi3N/XGq
pMNnIXqO1esB2WO3wEr5Wify10MWgG8S03GC8gmckjS/Lfq+6iYBRmqjK2SvtUuU
yRXcI094zvoTneyhSZxYR1vNhOW4Ti8Dq6wI+Zlj35GtTtF0iv3mt2dTCEDAXLBh
WwVIJFS1J48Riw8xRmVA3fdnSdECeymJFwY34uj5pz5ZAr95ZlFjmKJ0Hketskav
CvQIwXfaA6sIFyNNoqpgwUdwDsksU2as9lq1xU+xMAKUcT0Z0qDwK4M1krGM77LM
4BmWEMTWXqgmaEcTvOGA1onMbBz6lKlfZrb5FbuhBFgO8F11Ukm0MNT0w315cs73
jXKLgKznhsQWEab2er7S5SsjjFvOoS9k1voFvkMS3Z8V+BoNazJvka6xGO8uh1N4
6fPMNjQJsFv5WrN0tCaZw2QgpgvwMavwELWCSFdemqw8cL7NIaGDxzJGuVXFM1KM
d3HPWSG8hsG4yOZW5gzDguuTT3YpM4dpqp/0ZbhNcV5YpMOhJMg5Bm2/c9Rxvk7M
uXVForhYzNEH2/pmyIzPNyFJJLwSwAfZQFxZaTapOElO22J4TE7CWmdIeVmPcbA8
PTZ+ZTuQx5tFgCdDMzmsAlazDInhUhYBpDqGSz8Ibp2wJtkMzLzDhoA4Zw5Jawyx
8RJrCaOH38VKCVvmI54RKppckgA5X2idwShmD5p1UCbMG8W/h+GvxQJHoP4+PK0x
ZDhv1IrZEgjpKAK+vkPDZj+pMqkBdWzwH4Kw7HvbSWO68vem+kJhtZGWJdsguu2S
axmEs691/rwE7zhycqgvOQw6eCWoqLfZedi6f4xNRzeYsNrMl9nhOrWvL57UKM41
/sWuBGBjo5l3wiI3sWqekLokandlNWbGV3qR5QPvxVwvKClt7PevlunYytektALb
bFPPYnjFSIMUTEc70OugdSl3vi7vd8qGciaOTpu38z/PsWg0C39jrnFiLlbR0fUr
sQUxNPccQmQqSbynicfZlkroDJQ0BAIA0IObIwZ4wuACiUKekiofBU6L6pZuqHxB
xudKe1lLvMg0ETK75+Q0Cq9DC6gdMgRsKlQ6pj9mXzRRrdNGOM7KmJW323i07m4F
jU2pJwCrbX/j+TwBgTaA5doALX2ZwJfYjo2CWwKWRyUqjgt1+5ArWKacXBmYZ7ne
tpAxZlKelkSjaM0Hbcdi/BY8mfXStDeLNuEHNwDPrUngceFAx8J2MU7qRPMeXYny
K/srfuNtXBY18jt7EqTQAOsmxbpF4J4s5Uyq7EKzP9g/mDIeFBF7jxPBIgs+s0Zj
iPKlGqocZH3uQVB8/XyTApkjO+oxjTBLALlqbJRe2iaqI9gwxMjrSq4y8Q7gkhiP
PD2457qgvA8SEvy78p7s2x0pB4F4mNzOrFU3FUVLscw02Hj+aIpGKHfUKu5IcJbo
FSBZcRfJd0RaDYOhltY3NYcRjVFirCdh2+/XXQwzYbHDrxvb/NYEMQfPr0s2wUcr
Rj63DOBLelRyvwMjmywca8CJxtpNRUoV5+tJ3rDpiphFs7i6rBDbGmor8VA1bVMO
Uy9/6ct7Eu7rj9a6zXlOdfYOlINqwkmc/e/0x2vfABQtZwUBym4Q2ULqPd95/5ru
45gt5S2ivY+uS/WS0nqfgJZKXw63ndUXz2//7w3oNDEapYTq/e3KzuG+D2ofuQDZ
Jojot9CxfEsLs3vjVw92sFf3WhutkvLy2LCgd03DocopKiwy5wd+DARrr3n2sRpd
DO7g5oA7zP78ch7lXL7PyyCGj10yRx/e5XVyiPKncZfnKoU99RlfpnjjDDtpxV//
F9xj3BGJZs0LLnVTOcTDmfWC9rJfiuM66gU36dQxBVlMuHn9EednnQlu6NKcQmR3
b4/99SqVwgn/7sbXRFh/MAHPNp7H/2I5Q9L65xM+njQ4IWgiG9WTrge+MBl/GnqT
PXu+WjawGxIHyBvSrgt8OR8bXEgjmvp6B9DLv3GACwPmA4vAWaB+xC/aDyKTgvmZ
7OxGwbe7O/9QGtSbPa5Zx3XHZv18ootiGVmlKs+ca6hFGUF/ChddQ6kBp4rj/f6n
pCAnkFQ/MlR0ugSOOi2lYSnjy38selwtP7f2oQMf2vd/FvmW1oJvGElwVtjrhE52
NgJFrNoWh/qZoC1/F16pBg0vOnDP58qqsFJg7bpqpfMt0OkSwLyBVy/6ialrvddQ
XQBy6C0G68Vk+6fUvl34M3nfwxtg8ymqtxcbioin1cUwyAMiu8L6hXvrZfVPVIbn
VSypcMv9p4qtNlxrT+Hw/8fg6JGIv+rcULLKaKWZrzcNzZHCMrLLNU0yiUFdCf6Q
BYeAL/xJwlT4kKoobE483vOqG8jj8UPuQqFv1nV7906xTfV6vRuM++ZQ2YvaueiG
2A2t3Hlq3kRs0U6VxZ6axhCBBKA47HLSkCaIr+PXF8lh2SpClUjxOth/ntHhqenK
HyB0L+Jw7a/yv/MkyVjiW97wT9MQsJWxPRlhrUoTqFqL1AseJJht5KqHijo18lOJ
HG3moT660Nc/vWyvp6bFHxaV/WgF6DEPGU2QSDuiP2BJu1ysvB4AKkOVG6+NSYpv
pgSvJQ5LjS/IcM76Evg89/t9t24E7ymMYqu3OyP/LrnPnGjjDoM1W7PokQv1ZqpG
flaUsFmvCNVy2yORGfIKq7jCTFaGv36Cg5Uv915+wvxE0MNe+oQ0FmC+G7LAVJLx
MXiOCspqXNGf1YLv6G2xh48KUKDFNJtdejI4J0Eo6jIXVqURDYMIOye28i+BCgwB
aZzy0qrNla/MDNBLxbrD4UJlmpfSyS0CsNo7p4O/yN1lhB7nN7rFTMb00WgMQOqH
08E3mwTbJE3xfQllYljC/ayjJW7llyF3AsouIuS3LDuQz/jI4WYz9pB0/jKsweI9
HGWwUl2GJQXdvrpFgrNxcK1+DLRQdDce+1EwfEK94Ab7zx8gweChCbDrpZita3S8
Ulk4QCHb2oGDjRZQTxytuXsQ5nRLyYL5rmcB/eYdCFVkEX/XLLim4ywlT75jCpKP
h1RCCBrm7/05NCszw/0TJUSrTDggEudAJXPsePhXHarpOdZgo5ygOc6UbOzAoNhf
+pEbxYN3Vjbbiohe08yXvksHVup60zWx8q4bMVLyDhyhstCb/U5If6K55JheopY9
H+wrq37K+plUAC7cvRazS2EIbTMhxBiHj7gSWPd8n7k5e12Zo9fqZaE7VquosyBI
S2jb+WpDMZ6Zr1ECJw7140EZLr51yBa7oTIJL4fw3ZWYmtIsY9A6yHetoOizQuo8
xj5MBnw3NxId5JioIBXN9nFL25m16xPsjJo6HNX2BLOwWz7mlJdi57lvoykUl5Uy
ZVUHTwi9KZLe3bBJQIwbWTfge9nsIw7qhSfSLYFoPR6kf0ivI7JT83oa1YPY4inw
Z5gzt3ppzoLkoZVJ0oGvHHBH1hdotWscqeh7pnr2d2OnqeVwUYxxZKxvHHwzaWVl
YpOLJQm7yVWHIW9KvT6IBjaTIQ09tJZRs/KOGMe+Su6VNmTRf/pk6yL7QvzIw0IU
VLYBL5IFIqD1Fdi996KnKXGcw5hjZeyTsHvQUN4drw9mKUhYO9/4vUakrCSfsAi2
BxPZc5/07c4aU7Yr/Aj7QHKWyFAfX7l7uBWlXGGpnbR2dYk4BWXARXCco9YYbYUv
02yWeo0UU9/dQvkpCR5ETGzoRahx1zNxAvJ3pQuAa75JH/WW7PagVBWR2Dn39Mvc
0PC2GGvQio4mYzXggOQGJnwxk9F0RpIEL9wAymEcohc1Jt9PzitzG0QFzNkc10re
/dO20cvP7zQo9M8RPUpksa+bdyP7XEOwa/e2BWogQqZcaH5ueQbVU0TSc9lSMjtz
CAqThAEVQCGBuERr9Sih25n2cx9yh+29X7Gnweyvn/kYdoQiEDEBhUSqNHKMEEYY
zNizbAIGUgGNyjpv6eHOlFnr7AioMk8jRnBsTYaZp1708ONew96K6sEZZxCgT0Jq
0mRo7d9rlAKodo061USNqs4SKQBydVaFwgyvgr3QAICWeCdzwolgkGDY00YCZm15
1zlKImX7oY0VPb0VYpqB7XkId/a4TC5geqwHne6fARZx+B78/7ex9nI/c1oGwEY3
J/kaw5b6TWf9hntJf1gRnC5fWiUTM+IhqLgis6/WsXBB6a2Rsw0/JNuSOOEgxqM/
OlvDyj7LdWJCa17/mhjOw2AFZ4RguHXnVcjvBWqH5MUGGyojUPRe6PlinKrqwUzt
JrzBxq3ywhthYsFtcXzCjmenM21AL6lwOYOBoz5vl5n9/Ccr2Xxn1gb2ZIsGXGme
nii2IJ3KwVMl2aJbLkV13lGyecsSeb6FRuEljJW9STpwMWPSFACLw9S/yBFT+zK6
MZXFAmBbl0tDH9G69oEsr9XoOue0vTWTfLzRtjDaNnNuX4XUvEj4LFG7PubXd18s
QsO7dVgvoUDKqksb8hnyV5EE2suBw5g8k/efx2P8M7x9G/3Psk0jyWrYiZvHQhVn
3Lmobw15UVx7W3oT3oy+kNYlXLpWI5HYoSv081PsMVrD8TCNT8HT77Z1C7cINqrH
lo7lwNP6Y/eOjmMppfqUQ0pa5ymBY2/blBUG+O2CqpndMIRusNnTrF4vYKXHKeW4
fXv/d87KtJi4dw9fc3LvreZXm6WguKPNsMSYo/e1vq0Rfwt/Gy+PpNXn0u4Cgpze
nX4Dfj23oUuKtPWWZp8UJBjMl9dbKIyffQPmlUPqvvlsWpwCYY8RoMhoKcQHfji6
LnlMjR7PBTrI6hlWehJJAPwSvUohUbMVyQfLvjuKiDslzSgk5r6X7iqmRVlPv9VY
mRU5Hxzbz+4Ouu6Yj8x6hpm403ft//Xezvn0HaeN+gj4RlqZUa8oZTMwH3gUVfOu
F/ePRSMGcqCXssa5hYkWXSlkE2ZLXDNIPTlK0LPLiRIsm8CHJvyYj3UMbpGdZ7fi
g0ucORvr/0rNI/EaWNrzMpzbYgc8lqRorxUwKRR1tBFaCZM9LqDbm38gt+NO2PJF
JgCulWASuMTy9lmODz3LCV9HS7Rss+8Q+7igXtuWrsR9vjvXzpUtOggxyLXCaTdP
Ui3uN3ERZJUM+lDP8HytXAnRe39DrU/avhiLzOJsqhtUb7108PR2i565Kj9W4uqL
6YO06SsKLimm67SBAGusmztZB+9UL7Ru1YAMLmBx+pQ11Q72cz6+TgJftwpY8XJ9
0sXsoWNliY2gdfr7lDoDwPekltOfWV8et7TR18Iob7Ow6PumE0b5I+2RFN4qhcuh
SEMCAYKlK23+zcFczUed9nmV/8lbh4/vbgdOp+vhPCQzjf6uevugAy2TNHzms8Uk
3a6JC2aeVgCiDnEnUgwEQJP+V557b8oUJu0r0d8TObWuhLPBRPcxcVvGVqXnb5c9
je9JNRM+8VX7J4mirbhKfKWXnARvpj8ZgfLhcf2+Wj0CK8xQVNU61M0XPD8cz/YS
NOzNffo3GO/A/Vb+3Llh/SgErGEb7NBe4eCF4dUNSJyhhs5a/OliGXgIWOSfp8hL
qoMFALQ3XMerW9uiOsjdCL9JNqJ5jMtnOSURn/ZgWPXa7wgvRw1z17WY4qMzeu5Y
w4VTCrLXK4rKyRl1oIL/zWwahOg/2DZIFuldwmw8fMxtlsL7qBRsp6ESglVvlP5z
PivkFT3hospyAjjw4LoMrSDuVbwzXdS4FQTMJ2Z5R/ZSPp5GPfA92qrZjrHd5Sjb
PAKYU1y+3lrkOCZbUk1pZaoAnZDEDcANPDaIRExk011hfUs8jle+w+mdjwxrm/5b
tji279qyH6SkqSagd71d9zLpOLdMl1ahv8XCSOIwTsGVCx4mIiBtVRQOv0Jfq2h7
GemgJryU1gcHnqaa35xgPHnkZlvfzOp9xuQVRHv/MUNQ1qrWKrSA9RRlKrpmSPuq
60TmcBz4A4eOcyscH3MbmdkKV2OoiDD2TRYASt9o6sUFE+nLGnjBIUwu6oygTY2i
LAoVURZYkBftdH6Wnx/NmommbNHSSTHd9Ezjw9M9BnqkgN6W+Pbp6hmLEIauePB6
Cv50Z6dBBf3DcLHq/pIzN8Zv5Sd0DkhQ9jwFvST/YXD+fLTmFhaL6uPWRvaKP2cQ
w/lEk5bXDQWcHIAcECs+dwV7SgMPp960XCwON5/VRaWvLcWnfAqvtaeJtBVWxS0d
Sb5RnJfnQah1AmqMPWQpAWXApGag2Ic1pKYqskaVIY7S0YqNZkhRpVi5mCOVDsuM
CWEpkSBQodsPcDFC0BwpZ8Pb5Hl0G2ICQXOLDf9W2UvWTDtqcym/OfY79SrD/5/p
yF7qGSXyr7prYXUMf2BF5Y+aueQXJIlt5WnJYg5h0xZ/w/LvBicEp5hurSkiVmkQ
j1azv5GV6zr4fe7r20Qv5dsKUOE/Ls/9op5bhRHuItQZMxvVi9/gikR2yZqlqcD/
IPDpHzfq9uxhEUTOfgw4jeR8VPLrCIXv13jfej/MXZHCslg8MzaycjRjGu4X+8Up
A990dwyzZF3YsfZL23LigE2qvoerDEfrsLGo6CauQPtZGY87sFthwW3q1KmbmBwn
JM44uRcmqZUh9ZSDWgQlPUiENHbtw7cixVvfYTyyNGWuQ2DrX1q3QimXiDs/1DSb
30upap5lExwzlLTSVZxEfuaemZOEaJR3PxeC3dfenKnvb4Klr2cANksimVpZIzJn
Vhlf6CroCfIOGQg9lVyshDnxOgghViArn70jhjWn3lsQ7IWAu4CPWY2KP+MIAZNL
8q3sXaRb6w6TDkTYobxvwPy9jcvIpQUmhqBcZtM1jBQ5ZvK5hrJ+onJGJgsmL10D
QX0vxzMxxT3vqOyjy63o4ckH7DaMjqIzoOgZ2kkuVzuiZ1xlk2S6PhYIb2e6EAMG
zxneZj10H78L6VvuRI6z3c2ShW1k1cwRHZ4rQtMl7aNKFdPbSZiC1j5y4AGT/jcS
bD0FQ8EgLvB22kHeEcbbMnlnlc7zaSXdba1X+K58VKG3D7YzbTYSrJgaRUS4zovd
GxRCgRHkCREfsef4AZJrGuT9hwAjaUSWqbSK5ktqXs8qeX02yHsHaD8dC6knH6AV
8zA6BKCfaFdqcfESo9zsM/Nu8rDveVO1NNmIeeTDYQgI597C70CAdOoZoJ29cG7J
iefieRi3On9ei38/i8rl39HE1LsYYS6X1oVDiF9wLDAAex6m9dwz2Rati8iroabl
b1efdun5LR5kqjsNPbP0H1HjsoLF8P9KEknliEBWVqM0Bt7x5ybbnRV7BYe7xFDv
ZEP4RAa/hVUnl9451lZd97znbtT+x4qqRhCa/D9dH2KT4llv/0KhQ2P6h29pjZs0
MHF3aCCEMfH4JN5LZQbCC51xsU0BkZ91fscnMb9GU/REkskj0z2eXE+bGArKZ9H+
kyWnoSRms21YT9cPFo+mICncega9jr1FqtUvopnuWq/i/VIHr20PY9jKwumGFcJV
sQOVItdO3r8AQpxPGd5Et9Ulg4rysBCMCErvu2YdtDT73q7vCbKmGr8ylAjvpUs9
jFcytt7NCw4G1ZmVoMRO4yrn6PTPgdSWOiBSkis5bxENRx9ICXUwYsKchVrM8Lne
bzkI5dCe9+Us6ljniBegTDw9myqQY9JA4K8x2SWaC1Djo54GnHBSOXEM0PYCip3O
omgtoNXJD8iq16D/hED42BWza1s+WL2rCGI7flcUnWeDczHoHDFDMVWekJshQF3N
BPrnWZdI2i7vJI9+fonubDsF8u25a3wov5Gs2N1B/CZLL1NCcwriMOXjlgKr2odH
twkk0a2h/ukuAldbh5rWXcLnbJv4Hl4DGrDlPWqn2evgtwKvnSkUqMjZwWib+2fr
cPqvAKsCs5UY0ZhdmnnVwB1N7sFqqsBqBat4pE8PNSxRrR6vbwBpPhyLGcLTfKE2
PkOIUKu02MiJiggI5NYT4fUoXn335jh/xj0E8W3QJ6cXUp6uRHXLC7baV07ezVPc
QTMRXyqCTzjAZTLMi9p90aU0dndePHWogvWUS/aFK+8LYTm1fQrGoamLt7Q922JY
IBMNqt/sB1jh1u2QzP/OJQQ03Jk+nk6z9k2ErakD6loUHlRYZqK1lmQ1AjjQ9/BM
eHJqlKRbgIVJt5lcGAKdVZqzV9ObnndwCHBG4sKQELnJuaLUqfKDWUOml1LwSV0A
YF+Z8UE/FJc1Cxs+tTxrctlSmyEXlcsPBcb7H4yUgYWwOpKF57UOhnG2+at8eNqF
Iu7Yz+eC1zGlDoJHlVFmak/9ZPlNkz5xqF0O5zWREEsYNv+1Xni5Vk3WoohVLdJ7
w3pBpQMv9BTECRZh9nJInLd9UP0Z4RImUZr5NBEO76IZvDtqaFUo48ZBImkeex/y
GgB90MaXlIvejOEZKUw4QXqLEO0vi9NOL92iJNqN1lZ45Rq+uIEe0g/7CYnAHRmD
C8sruxpxOXqcfLVhjPM9e969yfEhnNXOz5LONcD1L6cJQLt6Ly1FSHU1dl8Rb/aP
4lXnOkol3Ik3VFeB1h8cpASeCzvbm9YYAc5fLOOqOKLyjLltIOOxvOciGVKK+HDK
/mMeR54Ul4viR6a0lcJjVUB8txHPQzR0GqSkGDx3abnUbRXFXh55g5piTwXgQUYQ
F7pygyuGkshbXCC+m8lf6Vl/nwS1PDzfBh4Tik0hoMzvQbOYwRAmmSsOERqQM7ON
O3eSElg7qP9nblRgtV0w7LJQjiQmA7TpxnjYwj5o2iYfeju6mweuDy0z+jG8SyGV
k/gGU1dgAnLH++IDwL9uj7iyFdPJYYTN5Mym/9GQJ21w24c4gvadZKRff/7TArly
r3pdj8iT9XYiz8LiP4IufkT/a88LHfFidU5e7gISkfcovClhBOiq8EgseEIis0CO
1j4UzEwRo3SiQxhztsbo7oWivPwnWJE81MT9HCxanb2ZoKlSTEteunQiUbEvWXVO
uyLtHKTXNQKzFwSNwL+f8G0Yr11DFACSJYG/iWvPvr83U2KUhewjoJUDsLwYcM/j
ttJStZAde7QvvZj7LFVElXirTH08AdcYXagYBfBIjlu5mNTIQD6FS2/LhpGP2Roc
zjkEqw6F6CP+7VkYfEtbLHWY25a4nVumQzt816mbkapmbukoh52krZ+xO+0Y+eSn
jk08D9JKk+1ZCSuAOPtOhZHg/11obkE507hq6/XpEuUnHqaDUpAwMRREnHywWrpm
rAuRem0Soa/K8vDM45Fimrq6QCQ2dCIH+d2w7ArXK033O/tprUIHAuqsWgFSC7Zh
B0tGIFd7YsuHQKULIN0fRw6mF4WKyZcl1emYdLcM2jhjrtCD8mBMlINfwImaVLBR
M4gK8rtA7ITC59+ACfbsbt54mWNQsjLSWWkadqibF8fS4jqz8eW1IxaXznjgRu8x
Q8sWecZrZ9LJhhgvquyP6UKLDXZbURMetgiPAw1Ly3lakzbf2NgSEyCLJXWaBXUJ
eunuLcfKqFK1+p+mhIkSSOkomo5dUbLimFRAZhRM+U/eWaYruKvQh+wmu0cELoGe
tDZE2UDEHLVPpDksHz0CYIrXBakTwwpmfwxLM+Hk4YVoi4P4vvgwEyS2uv08il1I
w6iUFci0xHKl63nkuzDVZAFenAYaDSIYXSvfNIMsllNKccvJDYfO7GbfPLZdMdEk
juhfM6v0GpZPve5CITL6uTWDHMJ/jZ8ygnD9SkLnSXCCXVMgMlp0QQRTrDrVVvZa
DkdzU6+kvNPqRQkEBegoP7aeqj2CDwU/JJhsM2KxB7cKlis3AOhlVOZIZnN8sYrd
UTYPYsAl5lWSAF13Oa4uIny6SZId46dd+gsKRdcIQpjjsucUX7LH9ZeGW/NQLnni
5/kUKI2ULf8MODJR8x/WNlnI+JZNZyWlGE2whsjCIGpEegZtGZrTkf5zf+DktdcY
atv1yxzZZ4xSOJbb1miNP4zE0GXW5kKVlFzGW8OpUtoFAVhqI5NloGuc+1+VD0ZV
e6nA1c58QbDzV5Ms1YpScqkFcDusZRUHfV4eI6VM2HtE32qzNDR1WShfUC9gj4/D
/hG7HuZbP556RJg39fanZMckmlrG7Kr0YksFNb0wGjyb7bgohOuoTE9DEzGGrDbv
DEqvwqGyndSoXfwlocM//v1yKTbTz+AG2V5jNzqnU13yrPsDyk8d+99DM4tZuZrH
fEJXJMyYgsTO/L5EGCpFsu8t4Y2Sr2h6NY7i/8mTk6r92mySoNhVNIQrqW5duGwe
VhnflBKdndoL5lqn/dlw/8cNNrEreN3mhvpeVwSGLSS161rmTa5PKHdmFbBU1PRm
cQcLa+gDuk7u7o/KatZwdPxVVtorPVuTJ2qtGIVaEsXhmQLoefWcY9eIQvA2L/np
Br7FlxcdLmroGF2iKwk/5NQS39/FEdYnknrw20DKQTr3u3s7ba03F5Oy+l+cQ+Ig
TGkgoHlcJbPx5p48WV1KkSUmTdpaF/Sx+YEsr52rWenGu8CEEz2Om6StKdDx1835
FjjlB87O2iwL1dTND4gVh3FzTvnmj7hxU0/44XEF5q7LUwMb4iox4y//dqYZOCza
qWQSHLwOkQaeP+DMddTHcfmjntA/MCY+uvIAxtZhX5UU3gqFvX7CQ+buNvZBimuV
qZ4eS9/L7RUGsDdOIjr8KCfAtNy9dQwVJ7vLC4eHekSBmD6DlIjPxgQSfUU5FWDO
WgAqEeta8wMI16669caz8kRUuF96b0PrzGxGnB1PDAPIMn6p/H7MplQUzUhiYm2H
dKliYMZilOMXCTE6COklnpXLI4EBD+zgGP9F5zyWt7gcy0IgtoPXTAWG75yuiIKY
wLdIOV0ew/QESqnnX+wfALWkU1TRDaWXuyQFA7HMJIEPsHx6DM+RkHGVg1u7S+Os
88OcJqh8e4oIPt44jGvAR/dhzuiRQfCFxXFkVDY3s2EMyXqPz58pnA9CcQXvF3Wf
nfV40BcMbviKrMtEZTPRAh7Q5BejSDRBWLYg9qO9tdyd4x2DQrt4O1D97Dzs9/9j
i7spC6rT3tSVMaL4Aye2hsnxeAROxXht+lcFFyt0tyDAytfpa2Xv6HhMCBRP5UQm
auNYerQlmRshmMzH/c9xFiVQ8sYGjsQQY+R9sHRDR++Z1wpxokM7NygWK+dpoSlE
n4A0WNBZB8mIMjUv+Oxd/DBQZBnVQeMxIZrK7p7Gv0FlA7jXE3BgA0KRqyxH+lLZ
qgjPHG7v7GG1KKU2QP7rT6fsIoxqmtM0IaMrTCdnPBvodLgEmT/fmygBb8/+pFhV
Q2PajUKtPwojKX/PmpgeMxNb8+YFjs2dJYPljgecAjpGtjWsdU8NgAdcsawof+h1
yks15Z1Ad/WBr3NinpxCjwFVP1emYpuDz8uUbHl1fe+AsFzX7/X5qKS+vq85L7n7
esmyt5CtmVhWXCdf8E0FEFT/7iPQOW9O3KUXsBIbAIIYrFYMTEUw+8p+OB9fm1G8
Wr7C8XTtCQ7E8Ux4U3Imts6182ME7STnP3SdTsoUCjV2WU9poy7waG76zaVA35nY
yJWFXMrqRlBy3PD0oJcFEF4lXq+oxgCh6FsqADIlwHkANDPBWOqeCrYrH0QYpN5U
9A71mwoDegPGu8gHI4wVTKzqh6W9R0pIgebONnB+3wU4RBt3S2fIE/orTnaa5Gbe
RtkQPKXavGJIqr34Q2Ots3c6gaey8rpuRpuXbWDIeQcUrGrbyMTOJeWrYOk/apCD
joyutc4fC24GXi1yLChk+QukAbWxEMWsxBMmgmm0eEHgYbHGLDtApouSm8IcO6RR
qe2IEnihiKI7RP3aWFfAZ+aNkJIJQFmQg4zTwQfAnftFVXXmyqC67zJln38us472
LyuiuGwa4iirOgiKaysIq7YQhlfhAAg5AbRrZ2nbcbSN7hKTSod4iNiD4Pw6Wdsq
Kb0kyFOqIuFrvOEZD72VDTc5wBisHLpRKwzgFPSvV2py6X2LmuauHqyZN7P9VJ+H
SxqQ2q//fz8cD38NqAHoHhTEP89R+vVriwmb2d5TQcgiX3xTkUggLBcmqug6dWVY
JA+mPZRrRYZzu3H/JcmzZZJl9q11Qz+IZcubrLEHYtinGXVm0IT0yxEI/kFhtZKp
pRQ/l1DZfKP4mYVjKuJaxsr5opsjhtOu84lvcxi2KE4rqj2DzY4cQoja2kAv/TwN
k2xX6q6PejQAwpgHlWQsxvVn2SP3Yk9ejVpveCW40sqg6SGyNv3Q4TaQti/bVcOb
UlIREzxcd38Ue7fpDrPRK46zw4kYYSAfZCcgx5vuGNismjrW/9zQeaRHNXW44HO/
IpZRJ3c+W+KOuA4QrvhHbOLpt/KvisxNY7hU3C+0u2rug/+Us1gl0kkirqWutNTR
B0xyCb+CjCEfQgGV4NV1re38Kep/bwBo3C3S53TOhdB+ediz0MwEZihof/fNR0Zh
GSSGx0C2ZR3gTEvPI7W7TNo/6u+F7Dkv/wjvc7AFlfq5aTg0BbQBkWa75YFu6kug
fC+miyoc60TrP2SYDIoGBmCIRR1Jw60uTtOYA9K7dprLFTH2oVJsJsR4tw9yJkQI
zzpnvhdNRh+8J0uOBynssFkLdAdmZo3IuYXa4GR1TIxzjRo4g+6OacU1+XRb+UYw
IzUw4Dyk4/AE+LCHy1uBLuVY9Hi5Nw6BXuiFcdQeaQuKtO4HR8ApzIdTTUPf7ib3
keiYOfptQG2eU4ytSz19tXDj7QnepbPpWIYuFZD+ibxPS4NLaTFNtgTpKVKGiG65
Wmu06WPfxVGRCoK3th2bid3LZpFaRKrd1jFjdhZ1nlD2T7WF7U1CX8yoikMFjuc/
KX0S0u9el1w+eTcWBVrps3KW9vJ3ngKODPLsDv+274GT2yE7tAKsA1BwggXSJHq4
ZjId62xcoWsPQKmZwUKzyChw3vJIfk01hHrKKviW2XdKGkVYox5g4gPN1RYaO2Ub
lq30OSv3D8bfhLrWDnLIIM1nJ18GUzy3ZJSU3KVHqHmQWpj2xaR9IdOjvgkBFSXy
wt5Qh4AhFugnixhi9mFaniVd4Q/Iqc+PzAGPtYITjqaaFXyuMbqrnWeCDi9Lp+w3
mJq+vqXLGhx/By1cqjhW/YPYHH35HNpGPm0bi6e005aoufWaKYRtgjB9pLcj27pu
CwPkRNPTwTFPQjQZtdcgACRhKp4S04DQzVlaQAevEJ+X+CfQTXDekKR6MhIfQtJW
aba/Nv3yMUlytEaepvrND4OUewLgKfbvwZEcG5jK7lpO4DZmEsKPBlwmXPjjfSIe
R9pU9wfRI0E9atBozJnEuH7j0qdEbQ27/f1JfssX4OA93XmKhAC+vz0MRhKKp7qL
jlstTFQ0hHpodjBWjZ+GeaYTjMAFKi091ijGliN8uSRItLNhDpBOtQ/3jgBm0BcX
ux01y3WEc78n9ITWu4/Rpfz6ciptStN2ONkBheGZoN5rU3N3Z1BbxAVLgrGDOy+4
qP/FxBZGM7xrI62JEuerVG2azPzCMbvKclZkm7auz+OPL29V+QYMlpA5XDYh5/qY
oACIRhwPSA7oYorP3y0MDOgvu8Y+9rrRVsMTznedGzFswNMp62iEo5uQ/rWHYtgM
qMUk17JHxVvEs9w7CB2QZpANd3pT72LSIGepGglAiviXWfeGvl4+F5CXNlxtX9qv
0I8V75q4jPvhgSyG9Hj5VrKaUL9uKW0DKGyq3AZgjxLAkmzn+PADzTx9CXdu/nTH
nPY4nwEJentCwUdAwcEtVdaAFoERij7vpavc+VHp9NHPnmdC3DIgs62A+WuSS74d
Wv5/2IZx25NqLf5oz43YJVON6Q0F20AaQ8Bp89xCnUWextQ6YBqEh6k/zVK4HSry
MTrgDxKTCYAdzMRN9KsgxCZ+1m6Kvsom/jFQpFWG67aoLLwCL/XC+68Ur/uEclP0
cm2+kZhoNGXbHCVDsTXUJWF6ai7N0fnqi4V5QvgfZW9Nq9T2lHlP8nHtK4f9qK+V
HFNB4+2YArt1z21rfcChlSal8zA9TpNJOs+QAyyqUPsXUCc113+6agnjwDK/abt2
O2eTA6pIZnjx7oJuLGBdIKSS0LPTdghK9+GFuN09aUbIWRuisv+2AcZxcMMPNxZq
JY20BlMNYSGbJNIu7uIZ3aVyBKdGjq/OCY8tbblTCOAjgvrGS+11Ck1G/1+FSyq3
uHAJe3VJhlxKHTDevNvd51H6BlpOFRMhr6s4YJOFxyq2ZLD5sXenX5wVkvOKW4h4
kKfKf/vVpXCDMJt7QqIasHl4NJbITv89XUhsg6dcMuGFrXeOwYP/G2TU7reyFlYO
oyFsvWrV1WYg+ZaFc4+Q4M9dLo/5wfiLfwQxXVjXIQ9hGk7wjcyO/qzkbopcnJBa
NkX44egJIy3dQlPG11dbWnHr4yTqjGgP4MT1o2HEKkdOtfuotJ77oWNZuZL6+ebQ
JdUwXEFkpnWCinND2qKweDkTvVV6amkXufZl4kT/sFGYcpU6PAR5Eh0muMJCfxbM
6K0RnkVnLwKAlI6bFHRujyx/u6JiLfsRRhP7Ni3c+8S9X+mJKmwCzQmZj7jpD2Vt
J/kfGMBSNkq+TaDc6HaPTgsGrxmMZim3PI5/2Nx+VvE992enf6qWkH3XHbHE/CH+
fXnKZcm1tKDh6XpQBRYPeNSoYLKe1dw5qeuxrSpanw9QFt1MvpfvMqfXbAyzPpsb
XQxsGiBZvRj/ggx9blXiYwdUT5Z0ABJcJtX122MoS00yZ7LFVBK1Ck9Lr9ytWEXa
IHwPdsbG0DyP6Sp8+tryb9a5hPiYauqIi1m1KV7uH8f78fdpKjoP7PNOSH9CUX/R
HtDVGWbcUHtxrInw6k6qCy7Bvot/F3cvWiNs3KAMLxaetAcNPUZiQ3lSG3legQd/
7RYPC0u/LcBy2vJLJLWVl0HUFZbeC0mzh+73H+iAy9Yva1mlFhOvw61SZXFxdO3P
/R+9Df6EnX99mxAwQJi2+2LMcp+AZJWFTwMOOEggs26jz4H09pNvIYxZnjVpd/La
lwwYhl8rGBZxZ2JEDb4tXqhp4GAE87J3a4D/RVWMj7FjX4veEmJ2MvaW5Rr0jxkN
zV76O7AvJxF3wVM1T4wWD7tMO+1aQA2HNvHSlMC3gdgEn5KXJ1zXZwsA3wlzM6sR
/KYitQWLKErtbYVPbTYc0SKEQbqDEfh0naiy2lK4nsTmUgfYFzAUe0K5C7xu5NiC
aREH0amwwfSnlTehY+LCjdx/cNGBQJ497UElF8dP26XFSbzti9TlWxAIAgGEYIL4
AgJR6oqe/B5jOXcpB/RcWWOHSA5iHjZ9IG63mtt/ZtG1e7SyF8qWJDY9WbXP7hYD
NOaY8zkEQnIli3MU0Q3I8KBG5HmEIC8tYtdfImQ+EbFGBR0FFp6+8jQccocD4azQ
0iqo+ezXTvCU8vfbsvk/4+o4koxKxalbkc+MODBTlxO2zkQcXXFhzUQOEytfhSN3
7ytbzdTy0Dq1uZVBxm/FLUE3/G5qpqOYRCDbRjy8t2HleUrS/xiHWTNvbwFY5+4+
rdu/JXCbqqrcTgZrErUzgjZMhGKIOfyFOW+JWEEDnTA/JMH2Fu1yGBtjpwrrGlb2
NE6lh6UTMXDEJHiuRSyhNQ7lafJaD5aSExhIzdYQ2lD4+B11ZytgYyfz2WspSR6S
Nj0gYU6EFKszsPaLK4ZNw94ow0BtcLf5FmnUFB/3Z6EiqU8o8yimnnBEK2ZEUNQj
8SF7SGzpggN0PUcfbV0OglUhip7T6hgMcePRnZMo4N4hUrHriRKDKI16S8mDjkWN
oM+WfvDj0MKsE7IznRHQWKfTKD3x3jrBCgrw2pYSgfg+ObUSMDkVOMD5EQYQZ6jN
D+0KXqLy4UFKZI6vDTppWcBHqj/bB8Iy3F0RuaTGeNk0n8Yg7uGtXWd80MFekG1H
IsqMHkp6PRWolLPkJKC5bKQyTKH0MJF4kKtQbJ/jbZEz9md3KSg9f3QMrshj73wH
pttGSghDpEmTHxcTtXyIhFFXWTFB+RWiOxZaqSlmIXtI8R3IR9F+Dyf1IssuR+9C
zBYBwb0p/14L6iBlKiDxoznHU0aHpxYYfjhVXNJVebpal5Ax5POeMv33lbUbA0g4
eL8bYB5oNQmI9OOQ2RtWi73BmLwMVv7wADoPLGHdFtgVxsWx8aRd+srlMGBfM4jP
tK8udID4CqxM46jFlRrwb3oJGWLHagLbvkZ0YaRotTPVW6UtsFcZZGhH4GGL/1QC
+IikmyA1jZPXl658qQK4lvRRYkpbRsmcBUTD5xrHj96W0q6D7TaM+y+voyPd0BdJ
z1uzy1fmhviAbeORdZuEPoAtkqcYATIg6HfrvLBNfAz9i1vcNZJzvEJAnk9n31mT
C9YN9h7OEPdCxOCbyBTVjoiPVipm+I589wR4zkJsRcWGyQYJWR3AOauU4XUmv0/+
1RxsDerX/a7boJ9MZ9uvQPU1AlxoLx5sLD+Zu5syQFMBDY6gaLtJkoiYqqz9XYUO
78Lf54QECtY8BmGu3pV+xjQ21TBs9NovVxzj0FA8sJAdYE1LNwxhDqCfnl0oPuoU
gXRYxviMBorxOnQICnPApPPKO1PtBUQUmazdPWJDfw3d7Zlu92djfM/Q2OWkXHcG
OnOqlsMOFwUf9DIomCvPvyqU3m/zbcyQIdvfMfjqkH8z4xhi3IKBO3H69h603hSW
TvKf71lx40v5KynSw9W6jr7/OY+TqQMgzgSe/p7P4M/LYDtK1G7iYXzQpxc+QO4l
4jnhwBxl48BjGRg4lZiiRD969g+QQMRZc99tzAMy8LSt5ibp7IWuav0AbVKPpaqU
++/mRoozoRN7ZOBWn1vY4VPhDeEG4EdGoiHSM/7Dz4ttaM4SkPAmc5PPdMAczT4K
22xnbJg6awaJ5L77xfFBKk8BshK0f1zq4ImTgpdWMsQt2vFkQarsVDmOvuMTUm7c
P+J9GPomBj2R49N+47LBmwz/lTWO0yJLBTpDAW1vqwSCjvziy9ADVO16MEwv10N6
Tu+EulfAgZwqFAA46lMq4sURkxYH4cSLzSjLPmIDiNe0tgzs9vFWl1/o8MNY3tiL
GAfRkm20UlDf6bYSA4dxdkPxUYyfUAqxvMwP8YFFjeEx04SajI/Yahw+ttPICV+K
pfO0l6jJPLNwbZTGdR+355w38zyvrPUnSvnVpW8L4xt16p+f7MMc3W7Z5gT7WBGy
Fl12bgnDLZQvWn1EIDmL9ZgP7wDLiihj2nXrlHaFY30V1LN3YRBFIVsxwucSMGwC
rY///IRLq+w7ShGUd1XxDLoEoCV4Guhh6xLmneL3tAjYIJ9Pgr/ZwObcv066LgHQ
J872EtTZ0Ay3+Feuy9GHxLcqYyVKxbTH+iqY1TiXa7JitjEHUO+sfjhvXXGu4QrR
+wuPPzYlZJYtt4KrSWEPCEQGfBAdOCR7wvDs1Ru0AxOF2EasYn1z17n3j4AnALxd
1D2oA0ZQQNqW/B4ksQdyK41mAhzqO1Ttqakc517iqEqd3m34pvCcHKVaHjmYHvlE
XyF4AZOX39VpDbOTNA/tiHvAeXMqvQTEVwaicNRwbQqiTgWWf2c2tTEUJ6L/KDXa
iQM5QowILhHQswKePkYeXlqLWPKKCHCRcOLUPeeatSeECCLj80bXiemf7fesVoea
ZGUyEAfekQBmdBh2GEHK6A+qgG1P0VhXATU200HtbCJ+tPLbuRar6g18I3ywbuCO
taqr9XoNJGyb8ORmDpzkDj25ARMEo+ejik6bOU9kTQDpksbO2vbscvUOtna9rFNZ
HFkuJ0nYDT6Qss29HLpvBL+U7JP5eOCyPbDVM/ebwYJgRxGJXOVcNkDZg4q/nUlc
qbCVIXmbCMwtB0U+Oc64mFTTGHGEUW9RSle+yUlRwYZp07HWF6F1tjm3lYdLGXYF
T7wuQmcUQ/l0YoR6OyK6hQ28yeNbK3m3pMyB4Lr0pvR/9yTOjDJPzvkO9zI+8BoL
NxdRu3X/QLVB61Qs5uUVJCMJYipGo1t39wnt4Zq7ln58RmYjBicKT/sEMT7gCeJQ
fJMWyScyDWbQ6v+Ok9i2zMsAgbDgU1Zw0rcQZsYY9eVwpm6l9DsG0ikI572vdKd0
0YWkBu3GBt97o/46q6tP6GLZaSfA5Vfn7vXt/MtUdhkUs7yc74n6HSyohKykRItV
acH8wp5eTve+r/Hp8a3Y3Z5yasqeGrntHJkwy9vD8dsmlMAircWkTCJShnGlasJg
RhuyisLQav6FRAYp0ilUkv46auMBFch1BssmCqXcQil2SEGGsJuqoDUmsKMu93r6
yNa4QqCJmatltqGlNLgNoB0Hvd5ch23YnUN1pptx07BIY5Pp0WuZIcKLt24HlvyX
YkQ+5DND0vCn6JYankiDSoWxRTIEMYmqc1Csx/9qFP4kWHdokos7v+HSAVy4i7dR
fdC+0TY3qgur2hX2kCJfO+SyAw5JHnvWMWbB7c4b6uF7dNzgQcmU+ZBjbK+83bW9
9wCJKPm/VnsEkbGfb3I5BJJ8r+mWlIyWgrxifNXfEEvYtMvMZuIgvGeYintYIXN/
blsThDv4yRpeYJQzxMJ8kVv/exLo9ZWxVh6G7PUBotH3z/Oukn7YnpeM40PGVHFf
+uP+gmFNmxiYSq077Onq9VmPWBrMcx62MqcYwSIOTpBVdmXSaupYCFDKiIN6vub4
df1tn75pzoyJRDtYmi6nq39LhNgY+YRnReJW43tN663wP84Notsujgo+HeIk4Jxw
ZWCeZ8FEO+KPvdM5url92uc6huMyLwpAAj/x2ci6n7ae/YtEmtcjML27J8Sk/zbi
CnSwm0K8MZKRHR+ZIoFuODCLJtFAjzkVQ6Yb7rkZ/59eQog6JD9W7kIfP1l6vKmO
Rbir2TaOTr6OQN8nuPGiVVMtKwMgDws5CdJXWJTBGEZZWZm/XzAOhjg47N1CDSiX
v8qvFZHtld0VdUDTyLxB71f1fITyM6xf5ufG5ewS52wkhITzgxj0qEmcgKqWm2BM
32qJeerQnxkZD/amfcHap9vFHn7SGvknvvni8uYntEB35SVHh5RoMwxK7GXb1Lic
uYb/BHCYuLxRzdOYQagJsH2Up3qLDGIHiv+ar9wizjXjYj9c5jKq9B72mtPZFHL+
tUKiI2okIz4eFYFVTLJrA9buR/PGv8NVCMGHaA6HPgBxFQf+DmFyewdTOEfB0cQQ
yqeyRBp2Qysq1bFdySZTmxJdMmm/zLPoW+ssDTzfv/MBHgB5tW3bClOqK3FPbeaR
Zu+psi66pLcSXVXJuxQJ8+9X5ZyjBfQ2kPOgqHO1J514u+MGLN5xWKtQrIDrqdVr
M65729ucJk0ULT583DNFId+c9w0jTuJ4iNpTKRr4P9/GhRJyRbAekYgd2rEn0fqY
9iLj9mnHKZT7TRPhreDQkD7l8vo/IxDw5T8GiYAOysBtgTyP4WXSw7YgOxOgBeml
vqkwV87gtn9lio2AU+R9wYhx48rDe2tDTP8Wndt4f6tvekHpMqeS7xXhb37PiXM5
jdh+yH/JRvCkexdQopLUhmV9BkD4QxzjRztmG/Be297wm6uuoP8dqRkizGNFt16x
LrUrSPvPzyvw2SM+TMw0aXuE0S/Fk5EeLieJTCLxnajJRORWs4bPeGQCISwPTsmd
ViD38D8Mb9GiASf70/MtaM6jHeYhrEfQF+ufvU+l2WqEV1IkSdkY5Nafss8spG+S
5zIZr2zewYy2QYCsTrJczqM//+COeX2MhuDrcXY3KLD2Bu3iCB28Wuir9aVc4WNy
n9uZTcuEBtTKdzo6DCUmNiuIFwtmN3ixGGdhgDv/E+n04C5oW6EQunR696nraLie
LsUqygAZQJPIcUTyy0uVLWZlZ6pZmduRa8W11FkV/4tLvkqfMb93LrNpIhvklifd
SJePn4Pan5ZDGkrXz5WRVB4YD7QDcLg/hptpae4ORdGH/YlGI/dsdx2YtyeNZNnQ
Xc/IUkyOBwOV2PQ7R46JACfHpOFOywdcPd6CatgFD04QB+Kcu8gIXg1PqvL9vFjw
MsZTg0k6fPowcat5XSqrctc1R3Uk6aG+c/6p+vZxu2j50y7GP0qFloYgH+kISDHA
lLaDmdFXKquHkCMRrR36DTFLTOiu4BTaQKTyx+/GQPynBvGo9hvcxjZqhAGQY+vJ
HqUVETjbqULpfXjTwn+X+0tmogctu6L6koVnosnsrljHTGcKXcjoezpd+dnovDV3
vDKCJww1ZcN61+EnvJ5MDD+dpn2I03QZMzunLVCkmDawaC0O7Uttpzpx6hYA5a3T
eCbi0oQ4OCoINkICAvQIHN6oMmd5clQxRd9e2gUoNDTMGv6YRz/Q8H8Gpwzk1vyV
fmhfWsaX2d9FxQBfOQt/r5w1XJacQXHclLZDIhE+edX7Q2fZYpCovupY4B28hnLf
mQlt1qwD6fuL+nxptHR3IVABgwRN3YbFLRb927sjh5499RM2bau4BzGdDMcNuHPi
tTHyo7Tc97PGwJk6ce8IinQW4hpox6rgxx+myuXWCoPQktj80/B9AzgnQfj4+kl2
npzJtPT5+ck+mWSOoPV9IZlNJSeu74K5RmIxl068m6HahQPyayjq3hwX3FI6HRD/
N93PASgjVky0JqXjx1eDqW9/ubmy/PCKeX6gmqNMu5Gq+cdGwlZ5BbpWQuOOVhtb
9BhqgFVD5VFqPoBUzaZQPQkctULsM01AY9RK+7RaLwIsInErJk4p0bCShEm5WA7y
7diibmWPRyxMvER835x4+60ZEkWwyheSjRsetp5bT9JUzS96SsWGKqU9i4ReDZO9
LylBJHrntQousVnYOpWxuP5MucREne9hR+F1RW63nPqh5l4bgZFr349ZgaVOtWBr
xKrtMt5UaBafL0dI222oTUxiRY6bexfRU29TCUyKBGQ46SmiY+0o1qkYwsRVAYmU
KDl9zKCCQUtMiEnCPEOwIrSb9op0z/T1ntfNVHh5Kx+mvF1mQqjl74bt19iPa3HI
IWhbAi71YSpt5K5pnK3TMfeQ0DxMVW2L1GQaOKNndjwAdnYhjM0uxQwsSruGlVMw
gB3iOSs4ytLIAOu7EDIv4p0tZvh2LtsHmXWVNkLYZ6JHqG8yMyWdYajPHBFroYlK
sHxucJiOlYYZlSDiV1JcXhLAbH2B1rmi1KVOks3OeFM7D8OMj+pIcrzgB7YHjJJA
wlTOWY1Y65QDxbybNsr5XX9IGAmgcCWOV+nWwcd00/0YgU6i/IozTfqvpe5Ko226
JyKlWeS60wWNMX//lwEeK+y2hboFEeyYGE7HZUhE93XiaztP+lMUy9NZscIi0iJD
hiVcQnEuz3YTOEdODl7YXBJ6SE/AeKKrdug6n2WN5OSKSVYzzXddYlwJQCtFCXYz
P93yQWt7JHSj4a3fDieH6WXsjBxO99AU1JBsCmq6aPyrPOYmMxekvvOQ2azYXDBO
ERu/RcXCE5/fZ2XjHQba4gXYS4rxt05fABnB+oTJGFxCka0cQ1+jyyUEvP0xRXa5
r11Pbx9MlSNGjkCRGaLGnFm0nbbpviVw/D1loPXRjSia9ryg6ZqduM4bG1G8Ejbq
6GjdzskHnTpmOX1SKMtnFTIf8ovVp5C/Ww8xKsbNebB2ro+2tcIoL3MYOhbL0725
h8vZazDnJ1oWfkK/lAQbPZ2kx5Pb/z/TMX5y9A3E+dctWjbElfWlGC7MbH11tp8a
Kv3hqqB5nfPcmb4Q34lz2RFvUxWq3RmvPeKX5gJcsyGN+nOy7HAPZ23H/Y7Nmo+N
KrPM5+PxsdIiVhMgB7tg6atYam3pajV7BA25mi4Bf6TPbuceD7n2zFmr1B/uvBP8
VMRzIvRu1DXTrdYzech38FDIZ63NVHU9EUxVi4zA7qvq5OS+StbYuhxxXgXJUL2V
9KuEdc8/ezIRPnFL8odTR9TIqcJsGkqGHCRRWpvRGDDS349XY5SfXtjP74UeXzYk
kGILC6utB0yflAuWEvTA1QPBfJptMo0n9iQVbZ/GCqxONQTAYG43zAEOHTC/pSyG
FxqrLFsar2HfSpTnB3+SbvaJgMgIuflQFC3vHsnu6Lfqn3U9w98PoqK8cQx1RU2T
bhVLqBDpViY4Vd2iNviUdnGK2NGBaNLrDrH6P+OULvi5kd35c3PucwcsB0T8fJKa
kQ7uGtFVYMQhxkUBmhJ8L2UoCnl3LsvbjP90rVBsTC4WNDc/IjDAS5R/lVQLn6uN
I+mcEpTsxAZ5/DSKC4iTqGpCMNfTHnKLWrgiwZFDWipZLftPP/sS7yr9K2WzmrdE
ST83ZM+RlB6d+U6ZVzjET/wteQYAIyNrAHtoEyRVkOfAbxmD/OX3xQloRQ0oyOpb
jsbAIuVpBDdWAes1dxYDgRkxWjZb7iWvbsHq11FEvUQhmx0bx/jTMf7bV1FE1Zxp
WxpxvE4TMJr+XCAM0f01hhjUhjxCCWBkkWT2j5XnXJ0zPKofZsbvCufvR9ZsaFk5
6H87r7HJ7/aRy4GuIBeOkfJ0rwkiARRY5N730e688/a4pp3/6ERL1DT3RxKtvstD
f4pBUIPAa3HU6Ds9854vknnhT/q0KUkaLG6HeUKGpHn60gxCye8Z88G046tNuUik
jEw+sZpgr1guCTdGj4Mj89jlsA6poM2C9M6X9mGtohQSEodrmhIPrJM3QTnIorJc
bMfUJ64jBmLI108U2NfvkZtVigVF2S9CHSOxQLW0ttVSxceidXRUDxPBQOksx3w3
AWDAyPfyZwvelxmlBwh9AZMdgjBT+q6pBf4I0xTKZGqMU1FIeVMZZ0j59/L8Mc0w
dqPVaeCVcRSCqNSqZn9T03Fv/bN2g/OOj+5qrA4GRDia5gzfKPCTvuvrBGIPT9+c
29HYwHJjqi4fGnfn2gTGV5t36x4rs2xXxxH0HU8SUjJPhjcP4QhxiIgN+eOdlXGq
tkfyadNH0ZK6Q7BvT5Pj+i458xC8CBZEAVs8f3lf0R2cI/dla11K/ShCnxR4K/No
PSPvhYC5/6ChsC1XfacafjF6OmtWwmchhKen6gH5o9IAY5v3+M7tgJ6v1kufLeGv
SGt9riZHQyMUpTC+SxGZ7VBUsMTNpsRbHqxJOcN+Gk4xNbcqU/55o2hZZIfN1zpB
N2fC+7s0q71MHWvrVGtjKhOthYWNFiZ8E4ptnkkOJKwGkjoBf6eFza7fKWyvCW0G
2M+YHvksyuaxqaB7t/jX6xax3Gt34bVxcrVhCNGZX0PzvZ4KQMRiryt7CWR4HonZ
f6C1rk5222xAcsHy1LfxTbFO+Oyo50EA5Juc665BS+9q/hAq9BhShpid1CE4Asl4
UV25VyyiICfpEpkGa1Ih9YVsRER7jql4s65w7OuqHJM5MW7fN99ZYRbwJQ8S4qAR
E/Y98xaL7oK5vRxTNlOSIGyx3LyPm1Ayw9M9UANgp9LU7RE28Q6ii0Yjga1URC7a
VQJxhu2Mrnk0tak/mflnn0ydRwDnh15UriGMDMXPyFTOj8jBHIr0jbQTnYBnYLtO
zpnDbG64JjYk7MsUdoe9mO2AOL34yZszIpzaWi3N+UDZRVWEub5OOkZjK64bXXjT
pduhJ6+WUzv+jbRsbosUCjoymoZB3JQuVD3Ik+H0/q1GAHI4phHwbTB9wULpjyR9
U0sUyY1MMZfkcdD4Z3RbsRv/akPaFRXn2LOFA3L1PjZiDGuYjYukFl/ekHzPjfI5
PR5prYNSnqJ4OwXAphkm9BYuSwSr+29y7w/bOMiE6ZjcdmSkE+i6ShNVHtKIKRRn
5WnmFqLOLd4ymShI64waN7j6jQoqrUL0xKHyZYmZ0l089Yh3MTH2af1ep0D1+anB
Q0m/O+qkdiyVapDUMohMD/iErN31pXrUd0UqMB/Puo0xJ2+a3kGqPg/uNE/YFQla
uC6oLtOGElzH+j/SmwK+7l7KO7p0v3h9OUtNKjHQSO3dcc0mSqYEVUWkGxacxDBX
/++2oeNOAbdsX4gudwn2+3sCBUo7nTMGdViQxnBQr09D57h1mgNvwcxucpmCgkJp
ZMJfY9m5Q/VblvyPgYPeEX6iR8HaA0eWhRR7R/kLYMeEQC7JeoY/v8x5r4g18iRu
xLELk5F35cYqZ5kSnGxsleYCob1gBn5hh+Ymo7gGqFqTrfst93Z4g2A/aSyp+c5u
A952A4S3uPK4hI8wAr/QfyLZY8mpco2fpXPyDqD/piQFgHXdHkVJbZ2SqppnBUMr
knjtV9IWKFzV3iY6DB+wzJVJPe9cXu9F9B5Y1Xw7Ws8DQIakDkr9ZyF7wGwrJo9q
NtqkJEaHSSnlbUho6abu9PdmPzXL0AM4cn0ujrPd9zD4RODZCDC2B37aRdOZ1l4A
EfiwTJzKPC4PmpmYTtc+CAKpK7QJTTSDWoR+FAOr3Xqi8b/oFsHdm/NGpKwdG21Q
j3tljQA4te0Csf+eLfMl1XeTFkv19fxgA33FJnt8RB0sbqSvnDZfLcC+MIbSYzWx
92qKTVB1dDQNYzfRSNvZzNJ8SrNdg3yyy69Uqhu91utqYubsyhmMabcrd3Yh+SI4
z52Ik+0RVfm/xx5O5rnE5FFSpN75jJDBxX0vfd5cS5bmxwbTk++p5M29BVCI6qYA
ap16i3w2SlBaq2e0Ar0oCzKdTTKWtYy3YIOJALA5eO6AOmF4uEi4vUmEWl/Z+L7w
wQepuQcfXXDJmAu08Hv05dZ7nzDQQkvBx7NW3ZQYB6ZjZRJfcVMoYI9V0xmnC1lj
IreaqHCnAw9kwc7AcprtDEYLXhgOv9xiFGJhiF6nSgI4TGm2vzNC1JacfThbz8/T
jV0U4PY4mfvOPtH+/Ug7l8pAPmGBzwdUDw7g1UjkCMxN/Qomi7IXRYJQLFrgFacx
eMPNrYe3iKs5acLrnYbGA7rN9pjhSb8KVzQA++rVX0hiD5IpXxVsAegfqzgtV9BF
WMqm3+3todXlUwWKVbNPy7+VvvgWBwTtU+qlB0zJd0GZ4hUzT0hPUgaCOp0SEs1w
EA8x5+xKzGcILJyHaRrbLkvgXkG7RSfX4xz/szyLJaTtzQPkBe4TmS8hKP7to0tV
Z8s6WE9tC6ENql7z35Zwz0aTUVC7y5txBQZoQnQK3WhL0pyT7do5X9Gd/CSzJ0MO
/TEZeYVHzgnNvmmcfmo/lgKG1L9OoZdEq6qbCIW5ey1UpF8Q65zvdKVSz7oNsy9D
xQ/GxzU96tpw1tJi+HCC4kmWD82xZh9FJtMB6LOxHQNWi75+Icqn0XiMMFpL1noK
VtsR/ylJdrFaB06OdpqdxTTQwV25+XQVzBpaSzV3A/+t4q2oQ665AfvpmP+ESxsR
afF9kQHRB7eHCjdrOP7QxA0OKcHWKObBL5Cu3Q6SWovTnTAkvFBJbbYFJzOS7cr7
PIw4giHmiOKWrr3kRQLGcVCjPXlYBLGtHfABPl3DOL8VHMHh1R/39XuGUv4a6I7E
CpjALwFHwSRwj73fckXcEwEnD1Wey1xE361nUQ8CzUjNm3wcTox81eTT3roqHSeu
xN2BgnpXYvs3ZTi97rOYdKlGu15+SkIz+nP6YDC8v3XlAXZTaHbT9vdh4O9X1jBn
yil07aM52DHdDiDDIV+aOILtIizcq/Oq6tN3rXzBsoStI5R63d4hop35UP7Azq6I
MxjmyK1fe34nrMm0XyP7WhBplvOdoiZxGXdEkiKyafvh/i5g6i3viXQur64WG3HC
iGFmVcvrSBCerR8Pr3FaoCX3sLAigDjQ4xD0vGxbncR82vwZzeg5HQssgIX0Ds3G
Ob7ff0b5iGFtOJHXliWnUcbbdHQV9TKozvngo/1qNFrPd7uC65xuO9AKphg5D0YO
fwR0kHTYZf6NNixVSn5wN8ElJ4Q5ec8Q8ZMEi/fDJ8C4Bqo/ytPtsVbVNURTsupQ
6Zp3z213BdkxeBJk4VtIDpEQTUrJ2F+nYlu16EXkXIQKtFETOL4wK7zZ4cu8USNS
ZDENy8QcETJtRWevE8PAClrtT62bxCzAI7lOWzxlp4xkR4oHDfYJinx7g2z+eOC+
UbD3JuZob7ELi8SEIMiw28W8QEPYb+fidwMRW5o8s7NvrpJZxps4N94BimYdJWBr
X8t2WM8XPtS6Hl7l5vCi0/3BAADsiKbQBxRIj57nn6WQLfXNk5PLVh9iDFr6w66k
oOahKESJwjL85naHKaMj2wOaV6D2oUfJzPK8quOzEmweuhpMZ3lrK8Z3yiKiseo8
aqFTmGLGKZ7Q3s3RRwa8ZBznIFzMR/0Qx0geT3ekRRIbnRgNrCwRkxEhYxW/xOJO
O2YjRl3lcMIPmmJlluZHJmgniEAukMgBC4Blbpw8s5QoANqfgMm/3ikhIYruzEfC
/nDERCHnMMK0cvtvS77abTLV2RjdIC5erotFfrccboo93UbfxB4mWoFykq28UikX
J2iXmOv73pqoD0VTyZCgvOBAvQoz2Vq0mRDZuNUaVvSODwp9mvTp4p+VCpCoYPlI
v4qlUgPs+0lcExUQxMQWhcWcURq6clz6rfXnQv+Hc4HyjT39apNdbbRkx04FsAkL
pNswVkIxnnj9u4YgGxyAAKKzxAtEZG7WApEPi0J7KsQLoLAcC+fUM7yzghK4p3Me
WXVS9sDTWT6l6p7DRQ/hENp5UG2MRDOCqGWmJTw2isBaEKYr+0rsAF2+rzeCXJ/v
xEdh4nps+p7XJYL0/Wkge8KjJ74+wNp2befo3x5wCEPWOebWcL8XQiUKAvoJRJXu
sr+6GV1CdQrDYc0H4LRynXWfwbq89JUoB3vQZGmmntAC45ghqG/KnSr0l9wKudEg
sFl8YR9r5rcl1RzVFEqrmAAbeyYIuo4t7fe/cSEjMgGA2WPqiV/JJ5phiJnADpu3
ZZ/SG3c9MvfzKaNK2fomKyPn1OQXhHvG6HCefU7EhuCKwznO5dACuBeCscOaIEcm
WgkPs5FL26XQkjr5MFRn3h9rwSqDhMdr1qRv8EK+0sE5MaYp9g0P1CqU3iZUfvOA
/kCz96t7DWmNpWUjxIG7uUap9j6Sp3Ae92E96wusA3AXzf6kQHkYrFFyjRx4M2c1
RxC87GCa8kBLmRNSIZUlL/SfmATQOFrPeIO0Bb7gt46stjnzD6+O2xAw7LaIZkvY
a6v0zQEX4AqwPFOTjUEPYU2MoQOdCcNVU6n+5YJStA8s2jxwCfzCbSPbFTrtn5rC
UufJGeh/zninQ5FdW0Flkz2fe1YoTti3R/CW8r7dleKx+WUO2zYPxj+Oob9nq6dT
90U10b96+TZwMqLCthc6/TR6qgrXkTTjtSypFglrUhsspWzYNyAPf03stHFAd4nd
zsvKsoio+k8yIJoHZSmgoFbCS2ei9b0WGyUjWlYxCCxT3JAIP+P25UzxQzYSQYbk
GsgnNarvY+aB5/4DlGCngG3/fB+YFWkYhVMEbw3leY8c/dma12IZJHTcHdT4CoJN
KEv8Hgvd6FIcRZcdroLoK0/mthCHa4Nv6aSbzjUJncXtWxRLMDLK4zP9OKEbQzFo
RrAIgkWZeTBgRNJaN76QZI7la3yC5oI5Zzv3LoSBNIYst0trv1Jl7V3gW0wSSo4g
bNqntruMSmBj9m6ntxtz+RUxP2ifbStYeNl3zHDb9+xCX2CLIoncdbzefkTlZGje
y9tEogEHkIqwNqT1EEzUr55y0OuAn6200WrxEKj4dQ0Z23IGw626SSWmf3bBPUJJ
2CjSxx1CtjpCfa/ZY58cb3YqE/avdgc0/R12nnYZStoDcAUL5FKIR1nb1PhDI/L1
jtBqLMxi3GNmMZa/ZuR+mzfTUmlSCdTajpktBndT2r91P3jUvze8y6EVnuB0m/dS
8+iksb/EJquX6w3AW9gO+MiK2US9OCk0Zbm6o2uHLN29uLl4pAbGXtiuzURcBLRC
a3RswY4LIFDuNCkkwHzsJtbTZK8KSuSuSCTOWe8F/WhvdW9libg7ilvNkY0mWhwb
Mvnn9QT/2LrBaX/+ulEPbXkpRKegTzgRG+RUz/XhdUNQJbAms2LerF7baXUlcoA8
hlNBxyC0e/G2/4qPPnqGPmf3qHXaygkkwBKW7dCXGEs8cTSLJkxSItZwdeNa3u0N
ALSDzFLUT2H8SG/2O3NwVbZ2rZTy6gaTBCn8Qfw+ijO/VL5BjM4uVbCoKTVfN/dM
DcII42mux/zYM8E4OtZjnYUGLplKGIV5p74lLMLEtOgBmDKLn7hJlyU7BLXVFgdL
xilE4a6hK6ZyvZx49nZfYTsOk6R0Zu7HxzC7A1rfp6mfGswGZFdZPAGuAA/6V7v7
eEsdYvrN6DcGOCYOwKmo7zOpqPE09pZdKaMUqtA2vMp5iIao/JwGgkjaJxlsS1+y
PiFi7drAOuUzBYitvULTuUG8mKqZUyvZJWgbA81SIgL3W6/VKk9gDZdcsTmzyhsM
P5hzAktR7fKBo8Nsuzl14pqIIDNj6AKodn7bvvIghzAqK5UVa2s7K1GdNUM7spWy
8Yg6MbHBxUVLQZw7CNqJLCTt+OPDJbZi8l/rqI5/w0N/3Edr4WYZ/aSiYlwoTC97
3jS4N0m6RNwbbAz90OBclvCw6oSu0HXWvYXXa+MOPxiw54E9uBUr84DTYxn5DI/v
SoBuzuL6n0i1bV4y7P08E52rz6DRwkiCWRlZOe55cw+kvIyWnoHE2CAelKqpP7sR
33ldbT9PCCFjF7X/MyYLiehZUn2waxuAxwvHtIDEezNIM+fdWdvJCSzuSavqyBUm
3x67Qh7ljnEIEWJTyZWFZ9qFmUA46nYHWl1Nb6JmCD0QCONn5NFVyM9hpYVbY2fp
05CZPNfAYjwn77qS5hNlzpX0oikNafk5GD81wV8OVYsJZytXQnzLYc1kJLS0MgjK
zB7HGHlwolRY1KUKSJN7VfAiO3cxsUjy2twixKX7tEvpBE2zjtiHdILZj2IO9a7u
M7JkDY36tZYKd4Rl2Qg32qdrzMXBsigYsSkUNwXPGwaXiK4rvOuPIzNvNacF5HPE
aRUCsUy+PRcE3XxoAk19+Q8J2ytMoPQubxuivBLxOMUhKN9eC9OkaEIFQgZL1qyu
ii5wj1WK18UPQ6ogMkz0i8E7BRFZBTf7/lViK9XaCcujxdGjBITLtFqj1H/gK0AI
bfu+VxwF17HS5RgGVkNXod8pvDrBp/OzS06Sgw9GYnPEdYxXMkyeWNCSusjEqbAg
Ht6f7xKAtpNOEqxmX4mgnzGUr4CBQwp0FzaP3OziH8XesALG81qkfyaPK1fUTx2D
EpnGsokF5cHAEIBtLRLbbmf2bUOOkaga/H+R7h0THqUJvHBqX8NPzFbU3ZSilnsa
k20XU8nvCEzxzerCrE+XjnlOHvExq2yzz9Vr2XXZuk4/ZXG+3f2aRJ0pHHFd8snE
tP7qchHK8W+Pi+XyvM3emjBV1g0TjLyePU8OF+qx5QJa5Th1LasAkXgxRc99fVN4
K7872PopiAf+Ko5pm59KnvBknDlpQCk56Y945osSj0KyOFP/8vM5gj3WnC2A+mXG
U2fJogprMQqPgzDjf1xFxaGWzqtdDLeLELguY3xQcQI8zDSmrePKhUVwP05habqL
F/FrGKVIgqakkMbfLUeVo7bKz2juElsqowv5TCElzEYeaohWK39Ieqh2cGWNWKBV
xb14K17Y+O3hWyUB3ZeI84nhOGDUHuJh9RA8JI4quqsa3jHdzwIldBTlIpn2ibhe
Hh/hPisf2VGlD7xpD8QEtoO6cYwFRODRS83GNrYB+N/uoT42xw0pI5rQQbDwwD7p
2Qp9XswlaKpYdHNUAxEqw/kEx9njsRtWOVHWO3YshxcJJ4GGLpKB81wyrgxZCARm
g4p+jfbt83vRVEnTtKTku4C3M5hfVWmKsfTskLTLsrTtD189SWmRhJXbtQxAr4JX
MkycsxjRziuEwp4nPCj2cpAERdkFwkzXsJOuEXqAiFcYh0GSdIwz0yDB2P/84AXL
fHWQ1fAGx92qW1RWQG+ioEQm9ICwVB3lxdlG4yyJIhX0/u7N/H9mfQ004Ik3k1L9
4hhMVq0pF5UPqZvsmXPS/P436EUlmZA1IsegtrN7scQLd22pUSko5kFqEJbva6LG
fZih02dGrr13LgNKQhPoRZSHhvbi4cGEwELuu5zGKyKqC4JMpPEKuH+p1hyma94t
+vnEO0j5XKacoM6pLgs8LWI2tDY50pLwoSDNGTAMF9xXa/jAC0o1ozJtXK6N/wwu
LV4Lsk40QwQS3xeC4aCwIMqEAFhROuhAjx0gHDXOQV5s9Odh3Kll0GHuNNd6R30K
C+1UBX/2rq1A8nuZ70Dk8I0Ioere1d+XQBO1fEmxBrf3sMX+nvvvUppEMvgPIHx4
i3Ze6F17bIZUx5gHWt69+2s3rgPEfVOmzVkCDUZNITVpATHH2ZGA3cZdr1eTSxBw
48XEwMWBb1Fws+OziRGkNeCDrgAU5vEIpZu97tdMHefW56shNd8Gt0UTyJQDRhj/
j2qz8iMeaMV+uCC+wywAw3AwY/n6ftx5Rax4hdKvCUkKOlgGAqohjI1c5oQF/Bfu
mAAVIp+mzZIxdAFfK5/rDLFe8mXoXkhDnszfUHvn+l/JHRM4FAEK+1UfdvNI3D7T
TiYbkCuP+cdIFfLgkd83hMUuZ7e/l7Q3aosW1zsBGQM6cDDBxR9c6jNPoG3eZGOu
D2rSB4/xqMJWLTTmwnTzgTwoW099ZLmzUWK1TklbnJcINqQ47pFgRaadre6qfcer
l4Y6XXCYmbhdYFrhTQfTimRsP2uluwGAp8Vcw3A7f2GdYgpNTPBUssiUmmz/Wkaw
+KKmKGbEpfLVekToE40uz7seJWXhWgfh3pGxs6UnWcoWVKMqDx8JQ1nrNnzL1d66
NwxZzliBmm95MIl8GsBROPLHZXRFAk6HYl/epLpo3Cv/AMqwyD1SMfjls+w1Ih1Z
vNHOLuvDMGqOXDiJ0V5Qfc7iezjwFoAmZ/RHbmKkGAX8qzdWqH97tMUb79RiUV4X
7Ah1OpJyffrqeLfzlVeISTZOu4/CpysZh9ssMY9zgTKxi0e5gpbo3UuqPDLraDKc
bmVZWjHEM3Hh54EkZMmn44rJDoUDXsqnw2F29NTDJe8LX0rITXJo6Y++nhvT59XF
YPDa3WZ3k4Yk/BhLH/Z0WVSpDNHjSYQWblZ8zd3b5yhm68l+P8DF3o/MI+9nLuPY
HhNhH9eIGr2trvBGH+br1ia4RbuVXPcKXCJlE8Z3JNpc4BiIwyqDxwa2SiGxD8M1
T8w/nOf4+ui+fOc8TuRJYlBvXmmc1woZvgk+lPmIoW5KyNkPuEqqQ+1Wqts6Jhrf
/Gu3jIpoFnbKH2wGoiSKLMJsDzV7452ddbAD/NHPEmZkqS6SiXUew8c4/pOAYOcP
wPsCRzWX/V3KI2XLLlHt6M5HLAq7tDc4lQrZ95KnzSkX9YnSu++l/ShPQIxcrwlE
y+bZAGushi8uVjxEBSMVtypDfifOlckiCTZZriUdzJmXUWe6VyIdAmIuWX82XWmf
YX1sdVe6q/43OCmAKRIno8y3bdZF9LO5ohBv9ymHWXJ2zQ5oLteJE3SqP9Kgmwbn
zeEB0hsERxOPqM2cnPEba3ptsGVBURsvlbbTSVrRwHOZgGJVS8RVXDTYnxEGbnMQ
3zM37IHhGRxkm2r+BDRhCzdRYTW+J1Qo4Fz/c0h0IuMYZRy9rWeZdFjwQD+el6bu
r4EvJuzwb/HQtKB0KUtCYsKgQVL/dxqHR/YhZmOWB1y3TEnQw3kjyRB6PU3DrDHT
AbX8R862sVvJ2Dvx7JInF7BSiJrXSP6/cx8siUyaSfRoNh6dWmt+p2ZkshsallFx
IItQxK7AmezsfDXA/yBtkUkBH3J4hdKe8PrpDw1XDn1GKi+EkUGF/2td+G2bADvw
zYGna2kHFZpduauHFTVuZpLwh77Yjsv6ileRyLCQugjBnJ/axNfiqvPyp8I0qvU5
C0I4H24B3zhsdEGiHfxudba3jOYWdG+ZGxPnn9QVTFvfmYxEiUmDuPpjxcCW4nBI
klVFBY6Ebff/pyr9xmzTzedPEM1Qoutg6Gjx8qBdo5rPQM4rT8JrqzzzD/Hbv3w9
Pq1wYWtjabL8bY71kfsD6WoI+vKbNY2LmsPielOTZScHetwIl/6R8+uCAilKlJG/
PDZheUUO8QkwYF8HUCKVLORXaMoTswRIP16jroviowtMfhGchHlbjMc9zAfZjtIj
6hNW/zn1LF27CjMxBPvf75Avza5PF9Dxz34iXNqxY/pY5KZqX1jtdAMiBc5PgTD1
B6iKEFBhPtweKZUVOemXmFCrGQYd9Wq/dNw0exXft3vPVzkK6og9LzAbH3eb2v+l
DrHk7W2+mc6TMasG2eqiV8tAKO/rN/rx0nseigQAojF/Ja3udgcU/N3+htFk2b6u
OQOYeKIjFUBxRiT0tVhz3tlMKDMU5ouZD+0BUQy8vCPz8vrmJtzOagVPCFd8zQTX
Kk9TIChwglKvgFtK28YAOUeWNLAw6u8dTTgbNfdLUN0xoANuBTlN6HhkDoHXxfOc
Advrq1TCzcEkPctjroKNIfd/sd+MbG2orcyI8rGM1XHW5IO002y6ABBrqj/QL2wp
sijGARuUNxnUni4evw6KVvGB/b0fUxoFzT6SZgPMV3k1mOu+4O1rlPUMO72iawrS
bXIj8rumoJAGo5B2ooeTAsBQnsVPGjzCuimWUELhn4VFCsnB1bh1KXbaYIS2qbg/
6ff0v1eWARESIU2rRV1GQ03hM1SIEWdWONhQ9mJlDajEZf33DDtD5ALEKim2MCjj
ipWVhQPsCmqOBOUyp5C7RmMovEyp4kbGE9RnDJjFT+jKOT4hddrhilQ6//BzpMtP
yG9i9OleXgGvJZGpuIsYG2C8c8VQsObF6n5o0T38xDR2hyqaJK3hg9kZzSAe3FN5
CPvKZN2uJ7WB985Gqs9GMsPyXjzXCH0VSSuaecmyWqJvHXsl4IDhaLPBI7STGVmr
9cM7BD2QONIC6IAxMj80ayocs7OfctidUoucKMWw1lW62ZnGJxpWppwM+ploTYpu
0/qS+Sf96G+bexWSLN5eKPdjYq79MuqP2tEOApKjwlacpv6xoqbU/DQNqzu70M4A
Fq6T7lzZZi+t8CwjOpt5pLxjEA1ka+f51ileh+CWZO9kyQHf3Jk+x2iwGKGa3Xui
2TRgMOqhUlLIxBAgpLGot516QbQgIsulNTYnap/KGu21LRB36NegkaUi/Cj+imKJ
rLNCTEh+xD6TXsVwUt69T30PxbTqEGH641jHEw5xMQhlbBsykBDpV8dvbXbp1iSS
HOvEvAfZVbbEb63rKwa1R6YXZRI80ySAux3FkwluxY+wxvj5fPKxBRhgPmkNTW6S
Oi3YmfCXKjmMuNwoNBFFVC8JNiu0Oe6xCVZIkuwff8D1ut3ratKm873sDzMebEVM
tJ1usUj7GKVUfZY3bVWFWFrHFxpua9j8vwK1K5kaZ95Syaoe+xOu4bRvW3SCOoAX
R8UOHEX030d39tiESUNJA/8YlIAtN2ruYfLMpard5vNHyZrwW5bu4JYvi73dIFi7
vMmmt6AUA7XILvAzy3L9I8/+Rx2T5tjAGq9koop0SFUWW0TwjZ3UOdrShNgrfi3p
xm7jbm4O5yIrybgWONfPmA+oc5aKhxEG9bst+/HAh3ps8LEgkrPqZDzHYufe8sgH
RXGlRV/eNdoZXjuPOI/ZZ0LE5gkWPbfiy904o9TwGhQmjF3YC8bJQq9dWf9xLERy
xAZN7QCK4PUtLR5XjoytoS2I2y5yVx8rxgPrKmAdsOsj+6ZaWZp++Qf9R5WMdOLj
8uPseFjmrmZYMD9iYf4LLgKP6dbiIlrjb82Dj3SAAWLGEZtvxSZtFGTs13SuYBLX
xWeNbMjmr9z+X7aSBLzgwCq9ryLOceRMTpf3CzzI0oMJmVf8etK1QBuWMxWJ9Bk2
BRLYLEj9gLxb54wwTcdq7tmamjwmMGQ/vPQtIWtT187PktfM11vsbINKDn18HAYE
3vRKFB3HFN99gNvgATusQwmPA21c8+KQ17X9S7JFBBVlDPFJKLZDHsvljAAFTybh
cvpYAcVLw/EUG1uEoxPWZ1ndciOnZEkRw7uF7O+t1EqzC6ti/V5bbl5e5FcwO2nm
PHPCVrrtdGFs8tCQ1jWdV387+sREyHkz0vs+B1SjUN7H7xrxDMcMXqtaZFzN6CAe
BFdNtBijUAPUsMIXW0GKtbRTSR934X2FHZxFZTaO43IJRIdW2qBMF+x4+QWLmGWt
bj30o0O5FmFNWG+qaMe4XpkxS6WanFr2L94GoRZortRFEdi/4je6Cg3KWCTEQVIq
d8I92X8mutbjRxKOxBsVz1719JrtQuvATxrM9hhcvF/iBn5EPEOnpPt+oPchiH3s
YE2e8Qkx8BJdi75PlGqjDBfMFeVyGCsiIW5tgABIiwtLvg0d0Jviyf21xI4//Tk4
i9jUwDZVhjNd8maFlQHvNUKrt0IN2ykKVBsH7KRlESjJFHw6yJz7St9mZZLrkh73
uLV8jzDhegKgrpFpZykzipRXgYkAd+29PM8QKK13K9G4VJtM1Q0oW0VQuZQU9ph1
FrvZ6enJtA1Xyba3+QwJVEOM1xspJozBvgsyHmoXmL+t5D0XVjH2+OSOSOyvNAYg
O2+SnyJEzy6/WiHoAbKnBlg0t9+ln7j5sdfSGkub9PfXoQi8+aukBb8AAMSNzlei
asb03dd3cpvESxjB0Y4KoHxltjxqtE2xykErCMfEJlXm/JkQSM0c4zEnI9Q/K9YX
QVG/cwetQP6ojtqrJwa20U9XoIyB6dDSEsU+hRsMHJH82uU0TjQgZPw08k5fr+qr
PtWpWX58xheU019gf1mgz7XHmV9PqzhIYDPfhEo/9axMp01M4gs/UpzfNzLu8oke
UBAdSbE1x3TqJ8h1i6lF8NHxhVJoRAlFCfv0XYqjuq2UKHrkgiSu2nMHX1K4yMbZ
SlQIrNfII1vWYjALBerfhpQLrDSF4B9wsNUDq1WAkadCgUhA/Prxa2pGsxZT1E5z
whMIdb0mc+JdPEuGCzldoYF4ys/c9DmGxtt9muXFRuaRWElqkhIsD16TqiEUsWc0
PhdL2dY7GH4kTbzdlJtJMcHRfjWE1yxfE4/yjCo9vJRHM3Bm47e7mnIi5kTfaGMl
jXr6H9SNXYNVybpbnw3I1Bz4VvmcbMfXVTKlbPUNCgtfPcaNw7S1XDxi4LkcKJ3e
caYU7TnW4XRpupJq/bqoOBwpiyY6ZhODaqpgGplb+KZSsfpZrQd6I4srD5zj7IkZ
sAxzGBfbKAHpmGPe0qZ4jHjM+4bcpBn3FKB6KFe7OyEIOOhg8+asIFYEsdd/i9GY
K5v75MTgRiwjceaIvVEXnVK1qK5PrleElbpQTwkq7RpgZ0Y4qAKprbvY0xeipJhD
+NqWF/STLYG0hZ4W3m+7gTl9g9IBgBrscFZ1ypu9nppVtX1dSBgnY1Ts9+hcUmUM
j7cUp7ILhq3SuyKGriVqnaL9mzao+IfwSYrTIEecJaKbMffxGbF6QPMRVgaXm+7L
BA2nSewq9Xaa6T/iIrDT648OR7ksVGCf2v6o335X5czUmkpMDEpzfipLK0yfcaMT
rgOd7DxAK3oV39bJhJ1jsJoLkR+v3EB3+iakkXkuZTho3CUKsUjkBDMj/xRZ7Xob
8YyPlQpgR8/kykJFXxsIOUMl+JBOxch8vOdUxX15iob9hFu+GBK6/su5+7VJQhjK
RPkMAsKB8/02yYjfdhpBmM1jDUn85rrQNuS1KgT41FiwieFymjHAI3W2bUClmIrH
/Z3D4hBAOSLXN01JfZi4eWt+NPHucVPjiWOpuI8+HPr2oDS5E+wIV3Vu1Kr7nTMO
+snU5OEvt0hzlagvAgM2zT/UCVL3rmEIm09oJH8T/XYgjv5YmibjavU2av6Sr0QR
eWRHPsw85qAQ1OJxOLLnfCHpp2k1e2lsqmPweyTnNtsjVKv6OmkvRwWwmU5+lCG7
w3IvTLOYJW86Ry31NO1S8/dYcsW+55JuXxgn/EXTzXup2d431U5E2T2rMg8wyhXd
o3GzdSKu6Ip/jQv0uaamkX1O+bkEgtztTyBxcWe5kiv7liEMzMm2t58WuFEE0zTr
gq/0BlMQws+ICfuoC+Mjp715rBjnEZ3yZyaMwBSXz2h+dzDSMA3kAsZc8no0Ow7Z
52nPsP0J2Os8Y/bywAM6e3zLWilSmha4bgENwx/YWYFlXiJkRUHftKVo6ZQQNwKA
HZ5OSPTub2o0A38bfQ6eAMcoyr44Tve6okjKjYOui3S2A/DGK/Btw3tliWP0Pnbm
5xUygSJrRfyH0EHHyRkH0ga76XH7WKs8L7aIOzZUvHT5jdBZyuVpcgOoe53PguIt
WDtq2fCUAFZxOF+vJKbVIVQ1aj0Xb2LzYpvarhMYyG6lujkOCzFPyGcmvO3VJfL9
4jqb2jk2XRplE1MnMquyxnQHXJf5iwbEtEJ2oEFl16Hfia5jUfJabvOPeCeReent
hLqBqZh7RVo73oa7IRI+lcH1VU7lH6Wa01lohiEyoOm20tCIS/WzRq+ngfBXMHew
fkzr05x7Sta9qx0dlwcXfjhnCc5B43uceXjYSMwQJ7ZDK1qlJ7sGfpqsx+KREcfy
Lz5cg9D/hebBQNKlJQIVrHFhuvJe3DJ6PPlSEyLrti1cb9Xaqvx7tBGsW2jLfUhQ
Uw3JbCbzJVJKUZMmxQOb9BWLh6aSlaC/pZo+ihLPD5GKfJwuor+elLpZeBzEOiUW
zQvqZoAQMKIy2DsIPuZwjIJiT4IzzWcSfAFojOVIUDl88qWOC2KfuhJS4AwnFZT5
fe1cze86McUxVypYD9DGV+fEf0NAYYOGELu0Hay3zDb+MkwX71ksQzIc/32U8fU3
Z/XxvYibCdXzaGHHxUC/oiwmJiLbfXe09qTeOrcfqJPnxThqoZrHIm1jenwpzSoc
qOXQAmJd2qdc3aFWPKAIZEkfw4fRifOtNwfVjNeFEC+D9PV8KtCna9BjQdJ6HfLB
QUSRhU0Q0tF1gqn+HsNLKrhokBlh0YiDr3YrJsNfJZuH15xxP0QnLI83WfmJPM8b
Jk0nt0IdQxZ1tYqF+1nEuKeEGDxCLj2CcqzdAx36PgEqbOw4fSPqSczkKPHavCl+
/K5meHFHigoD+quDCGzjk97Mr7C1mH0+CQR3/r1cP/nnEQL3WDV4u0cwvw8n9pVs
y/KmE75l0CjTUuLzZDk3bma+x6+CZESTdXCpt6fE/JGgSfuLpOmdlnqYO3joiBKf
G4QpOdRHGBTt+nNta7b8fhNh2O56jofzp3lL7zR9QAXbilRFyYe7VsHo5Q5/el7J
gjXOmF+xvy9Sefc+fMM8kl4vhmkstl7FQ3N1Rf8E8ERDW8wTACDjvu3NxgKemJda
8vIqVmG/hlAo4gMKDXKamHe+x9Bj1E/vyvijLA1fkAFFpvYTqn+l9WhEZAJd1CxP
CheQ5QAwuWrZmDBNpAwcbm/2xJoscSI1pXZj0/tgZ442rv561gJT3UjQl2B/7t/1
IhmHtqXogP9OGAWDsk+Ym/41MiO3t+BuSc1dB7/YH5YLDuV3O5QYIg6GhrXs7kQi
DJ3+pCu85a2bfUvPIEH7ZoDR+rRpKpsHCUbPaevSP2fxbwIVYYojwAC3Kcw5m0yV
+xzITqiRwEL9bqcHT6IxQvxPBxVvOjPgBl227sRBG+vl5ruoD2HNIAb7s063CczO
3JgtAoXdaui/b+bUMfkluoNPJvj3tKmo2EoSWeWe9mkKfE8Ou562X4Fd6Mb+p+Ui
wnhZyw6P17cMkRQhov+fU0xEB4vFvzKStX+psbDlqmsR+qkQCjrr78hqDmAcc+nS
9geP9Y8vPGcEM56EYhkf63kckgqWyQBUYJpSE8ZQr7gBgY2vf5PI4cMCdANfWx5J
XSJe0IsfLQKcYBC4y1fFR23n0S22r8bCbJggfKZtXgI9g7Sy1jtegWrbM8sbQVjb
+/+tylr0AvEr88NmqS7sKESYX4mpYnyMywlodLn/VxsYU8XkG9UgXWPYObYrBkir
vTosBsgmwMmraG3YCGLVFG7OxEp9uZQXfHKxblV5Do4sXNQVhwNF/Co1CKdFjx73
f4Q/GP5CqrS77PVTWHk6w4olC/AFfradrMf+F3EQ5OImEQ13u2r22N2hUm7gGnkN
qYWAwr0NlRJAW29Bu6chC/VzdcwFE7QuPzJ0SHgCHpwrPwBq7EI4rWBLrRedjVZ5
Bld9J7cE6ZQFnOcaebR0aZthu9UHi+U/afxk6iAQswoVzxvItMV69nXuivnwU7n/
cSOWF72RKuEPTaCwf6DvoNhL2PCdddfj1nFks7EVl3XkhFXWseiqWCC2NIeqC0RO
AhvttoWZDaoX4DpzDbchS2Y4+JbzWjMmkU4EvRqkNGMwiiGLRMifjJISTLywPW6N
xfeqnwAy4VyIBi+4MkOcXhlWcoD7+E/PoZ66umty0ZXUDL759UDvca8aVpMBjoox
yveNLMF6ve2spXBhsm+lMEiCb6kP1zrRraWYmL5htxOy4qEeWqAMHF2rO87L83/s
M4AxPIdrSqqWYPtqaNPUHwBJ6S517WXSAwYR15y3X8mX9yIoBXeJUuW+W3F6AILZ
hLgZ/LqP8NDhkjICebDr9HVNeMOtTekV23yeiPVeSjYW+Ajqw3UqZxzpSK1krGJw
3yjJ5bFnSjacll1aRdMRDegtoaDI+bV06reps6w0w/DVai5upx7QkbYPH1uWTvZV
H6LZDvvShrfGZ9HxtRKDSU5NlxUzgAX/J/K63qNSqSvugtE9JMNDi6+4SlvRaT6b
accx2Vfls4UBvzC+yINlDiJm47XOLqbuAajYwNET+lpfwpS2muq0DEftXEZVTuDK
jMgkz7vXJpZlmYr3SOZL05Ai+i0zCCXZ6y0XH5kgC75QQ93VpiLeGJ630T+6NVot
BPhTP6vQ1iIbpVjCLWMkSvHx23DVogzKamgpjhBjVieTHwL7UT7oNvxnLmBgHszJ
AEUjw7PmLCrkN4SG38E15+nBsnOZSiqoX9yFyvUm38m6p1Xym5LNjMOtTTFJvSVe
JBtnnm7qG0WaIpqswxwlrg+c4/Voz2KxJvhUU32TMArFa9s1SchNoXXAiubB6D1+
dZa+IIJv05Gxh1Aj7viXmfRnD6FjZjsCf/Wq1oG8dEQAnZZ/JU9zioM/+d91RJ3l
PpaWvPBgSqwpUQU+5cTdtD0pV6BRNmMP0V4LCpEGqm8L1Nb1l5N6vYNV45LAFcbf
Km+m4TsDvPFQ9QvqD9xJMbfN1SKgy6dOwSXIF/rLlR3Rb9PyPFOuAphnabyORipr
erSKk5mmJAgDrgiglMSARikLp8o5SaOFFqeAT9x8ZTv75EVFfIuIfaDUT3NXNtlT
p7icO3lAhqHJR/NO8UoDKLmqqQ6PEzktPFI6Y6XdoD6fA+MlqklMUcmyB7CTo4S5
8Xan11/StChls7zbF80AiyzbYSx9E9HimntDdPQlWe/W70skdmN4pmQoxvks/qKl
frM+L+OdBC0Tp+LKsbTNn+Ve8466k+CyKj5lVqV7us7G593dlMuH7asOmDlNzegr
gnT1dmIyXg0ehq8AwDxDae5bwNeDQ5cVVI+oRr3rubey15TBOiVL1Tm1Dp1f9DKV
6y6b1Ad31GSX6XCFTVo1w/SB8q49SIXPx3FmHp0L1tiSPVNyyT1LIIVPQ8M3ZlFz
xyplKkGWle+tCuOEFDrsEbY07ZoR0QRzc+lD2BlvTpepGKns1L67iNWCKjEP5qYi
T7ZvX4y8cdt/K0g0ffcKfwN1W/0OtJQSCN4iIqm4IgiPhLk51SISpcgF0yWHpKu7
1KL7MdsmWdJWkrTi83xN/BmTsnBdlLrAOfA0Ao8RV8tHJLkdbVFqO4iLdvrKULnl
lzTXHcr60EExytwxYoGFxYq4QaOVwY/UAO4Wt9EQuncGseV+ggIviJzm1rMkIQMK
WDVm7aWEgHLeYOWqoSAeN0GdL8l/z7lqf9pFY1KDGFLEmYx1P0UKrWGdEEMopquJ
nuFSDKzLtPHVPk0F6IyaWY/nPOu2n6teLrQ1Tgyd0Iy8cYKHEvrrlNzpVehceJCb
S1xp93V+Y2R6fWl/8gLSfIj2Xqh/2VrFK3iVy7UqNfzma8FFH6nmE66nCiG2kdoe
Fug6xbsliIiY5UNvOCIDOX4ya9gToZ4LLiK2gWdj0nzF72Eo9HW5v3xnfw+I2VOD
1819hxAv4Xv1PR46AX9RzBQVFya7XPlEAxfsJiZPc+5xhkUqFPOGW8Z6oyVL5KYa
XIEh18UzAA2Nm4yBe5T7uNmb+syUo7UTtltCV0T44jjlS/NHypDmCjsZb2uAXfVH
LpxRmdmTK7xNN+JQT/R7GYBzd0ahPe9ijBNiW1ihr+ajSIVAO2saUmUoCq0fMSqu
bxo1x8JSLM10K+FXvQsDQxCpYtnARnUxZ87AYmknxBecPfxciNxO6YFpMbiEGRdS
eAqokzX3O2v/ioYw8JHdnKqelDM8aqYrpFJ+4054itKvME7WMa7UQnHIxw+bMygb
qimRXjcLjqkvyc8fJcYP9JAg/FW+K7A89UgWglE7KD54o383AlnCSLXarznMceC3
tvioYIz2mNapZVVq266rbIvEmSEBlV+U3y0Se7GVZ3PE2ATW0idfBi2RmtgvON7Y
jXqquyx1M/VQMDxd7mlAgQoM68EqEVgPjSzA8nmqKzVGpC7BKf1XEN2gAq9gn9mN
z0EvPc+6NtId4mO/d+fUwQ8b8jdRChEpbaMlWX56gKrroEFgudlPqXkgIFZbZr5i
b7KggzZMD4ef9CwSQqHOud1zhvCpE/oYeUfRUflO4j80u4YRFRiRd5SgOb1SBwp0
LzXosNCZgco13z6lmcTEBd9nixuqPel2ljupWmZZR4K3S1muuLx9Yypp7zDvzu2n
SSjXRc1reMk8ci4rWolrPqznAo3avkYVRWKLTXJGUDJSjEiHzVli4Dp0CCk1HZHH
BSCMpPibumRKPKqB/Oz4mO1nRre38BRSrsq8AYaiferthTZqNJ6qVXPbSBfSpJHI
dCABgR1WUIWDQasfaVmYKPZJ7Hscpd145bVpxmzcz3OZ22H0CujFZD+TQsCGi6P1
8OgmSY/C7MWL7NJvA6DTh5sKUR98Hoqj9yrV4CjQ4AcAJeSM1iVakU+QhSgN7dkM
Oo0sLHZj0YWkocq4jn/8UYs++Bz3LmNeGjzjFEpLvq9bjsRKJe9m7d30eVZv8Rv8
seMoZ3RmKN753elq86UJML4if8Dd03ihKBnjWmJDpdbFWACyf3OmYG5MQ3B2hl74
Ds7cnZKbSw6HRkOZNbNrHQdM5p2dnUdOHdgm5QwNEZoMX7xg6zLYhjcmAsEs2i2y
lKEpxXH/iP5Fe5BURu4iWf4bYUr6JZDVpzQtaWMP6lKwXzUg0D/YzOr8kxm7RTvE
8/sZ1AbRP85xYuMWwv0bB/Os7y/i3Eoe6nJN55E7BhAb3+uBtMB7cHCq4Y8IOK3g
losJNNyrRIqEo6IVdM2BZyJFJJ+6G99rPMdqIu26swFBlDlTV8qMPfE43jmjHxr0
Bp3AGCrK8PQS1baW8OTBDZDQ92RGPu+4TtodZO7lA1sfPS92x8o4BPJH2wTw+jZC
2+G6wZT5q7OIUb8G0EQYtdVk6unUYmnsq7wn6djJEoyrOBn1IriPCLkdEKp1VjEv
DmcpOR+gO3HUSm0/FQ3hkRWoOLuWa19ftVqKIbUVfl8qHAs6jvE/vwPYJikpfWEe
g/xEUgZdrDxHgG/CDX7UV1T8RmtfuzAA0Tr649s8XXSiT58ocKNZMQ+WtIYaZ6Y8
5hAiKaeOAUIexMDVHtpMXPArK4PHgBZo66JzNFJwLWDfP1f6ZbAC+OXpIYM1gOTE
GK/Ysk95eIGln6a0r20ZEvgGGxTlqbGDKBU3X6gxbjXve6Y8tbh0SnKTg4ZaCWeo
KZPKLVeiozU8+FVtS84hrv9FP+1s2eAJZzM24LcCuhY2+g/1wpzP9zP1xbBM6xPS
9S/llxjlB65Mcn52znH/ZF5ztJdhvNipygg2bF6OTOHMyZIi826lJW/BTMHd6vT8
Ndm1T3uwDZi+nFt/dBzspOav3rxNkL4Ew9CXZHWRiSRcDeHETrNUsG+DPkoo1/dT
+QM8nIlgHmWiDYHiN1mWhChN5YyzkjKfuHnIuqI0i9DTy0nR+hqxldZcRdyUFIp1
1NDVGxvhaqhhtM5bsk+Dcdna580bvLZVmwN4xxhA22SNIpcsafdCyAaXnRpa/J6R
1YWQXMjHSvmiRDDkVo5aAvhtMsmEQp2wPKzmsSzsDbJKY0qOZhbJV5mK9i+1p4zD
Iep+q4k2l5957F3dKknLpeE6V8gAs1mm3YcQA9b/rE2a0N/mbLzFL4Thrul7szBV
qqcPvQeLh2kydqsXXTGN/3eJH3Ny4r32YZuT/dELT84RKof5CQj7rnW5iFBxOwIE
4KZeftin4eq+/iBBlhKW/K1OCQ5d017lMPgzTXq5s5PUGhZRvDY1/dqet3CWErUz
byn0qsyZQkoZvk4TREtQs59KOJM4BnXUDdCR3h49X+ufHagFRFjO8BdD/83i5ysc
L4j+bUzO5r+kPnfEnSyJuNf+7PskHsDoKKUVoeCoOve8HBEsqmUghYManSv99pBA
Y/7DErYkTHWjwQX0f4MRkZ0xJ3KmVSpdZWSDubM7Xafr+JiFcC4AO3cHjJ1pLzFU
jRxg5ZS6EJEuQ7uyspUBfhuPQqx0PciBKtv8/WeuYo5Avy/fkCxlk+SdWd0bhWTJ
LHfm+/5pqB6s756b8doZIAT6c6BuXWTLoMQOq+yxTq2olBG5GCkyqkvbtJFmVCpY
OewCgbBxOmlsPcCFVDcfwIvzJad8fGa5Gs3HmZmnbedyNCjQe7l7fw6jTVGP8mD4
sBOZcTWC/HYBRe29uRAOy7XkP4um3FEwsFCeMA10j/MFNWowjuTMizKRSGZRzoj4
coDUXg1sitizyhJkUep72Fh0hGknMeiAQ+KtQHLJ4ZerXoZP11aA/pIafx7rJ36T
3amulgqjQ/KzdPIyFplD2/yaVs7cAfCqF0qtvFXLR5E7wmP4xp7//PihSIRoI3F+
b4kqbKsbiLqbJ2wWXwdljd+x+ie56EcD6oe0wz339mXswxT7n0E33FmnyiGxpq/1
Yvln6LtE3q3ASfgQkj+7ggG/dYPTXHfcB2nyLhPKhCkPXPMaNjRFpN6zhFbbgb34
EjQr7QG1/bnX6671pPvYs6wNNJP842YfwU8RjwDPljskWTXe1AQnAwlqXXXhCzwv
7BbjGiEqAtUhJFbuF1H8fw1dvmCXxGsNjQLAtLXPugvfox5tT8QYz4qp9LbfvsZ6
kN71eNjTZ8HEk4u+xXvFjcXDHq/RvRvA4wYgPgpWKgSyeeZbPxIpK278TWN+Y0Zp
33YEkqXyi7GaFP+diLjBOUwGwOFMqhsEbB/uwzmByq7wSbDgB2yg+fLB4WMppJK3
/SE3mmFgZwC/13mj7PBJPK9clTjM2KoLuKAhChKg6/TtdNXK+lhz+5Wh6I3H/oh1
O5WqNMP4jvcImyTerBMWPTSNX798g03P7mQWDoOlk0uEbxY8QV3nHBtxbmf6PE7s
KIIeHVrqADe3H4uk1DP3qvdiBIkMtNAVTiLzB1NSS35ScJ1F5A20HGzPahKkdG75
A9kvWRRXAENs61+M+8j9laylhNtEeHzLS/Cb60DFeRek7sfRJu5SNIY8YROlewK/
XxT2NjAC1WaZl5qct8+bsC8fFTr0qor4ioKcT7O5JVI25WfPK7oZQ7bFwJAK7mq/
wdR+fns0PB4Qx2U7PFBvNAX8pcf2uyCTBrgSMZoMeKOgBTKoWEP6m43m6QVLg4xR
P+9UpcaqaEZFg8yvBd5R+TdwwoaI5H712RBbiU9le/knNo0531wZShSZeaxyFL4/
PYV6McLGZH4ECFve9gAJ5lpI+w8a5K09ZksHFNOMSylWPUxYNhwpmVxAl926wgal
OD4j00PGsfW2cRwIqg6RE6AxYRG3Gu2LJkm4v6XilhNgNvivxJURFPLSjGs4dF4j
acd4tQkzoQc6Q6MLy4qgPAD0UJKW8ofevT5bvwCK/0OkGksdr3FWDrFsQg4JptHT
u65hQimoWgXDL7IGxhYnb/TNjFyUix9g9cJj5WGEAxXSLd7nsJAba+5LP51NVTYu
YXlK8PSDatpJ839yatVh+2lKoj0CeiJLEOmCU2gSmTGVmnIRs0Y7I33QTKkJBYEO
/Myp2a1LGGEpzvSSmeNERUJHbUKK0UvfV9Pwcg9DHhmFSJsaWW5EbrUF4jy2ezXu
G+XEt2SuDyrYLwCpdHxdXwkX5HpwKN+faR4h5XAHTA+zp5FyvwcapMyMwrgO8Rs0
pYblh/ziT3V1cyp33/hOmOKFo9sXx6T9RcjyzbXarDj+7tTKI62RrOEpsUQSZG3U
6i7HID3B4hRu/Dod9FBAuO/uNu5jMFSq7+6JxXcwlAd72b0DEFKwhQ1TX8AE1x/I
eaZo5OXlK6890m/q6hNFJw54p+WwkY/IufuHCDdtEIgorGEAaGDNFZ+MusAwcEuH
7Zuxfhai2EnGJ0sHZzUlsGhFZdxt0JoI90LE1XEZDDvVlkkP9LHr820HnueGT2xR
XYN+apsglehX36/pQqN7J4WmZFWtEaprlSKzmXHK1CTa8kyFfwGr1p6mWZ49jsEg
3NgdnuKANjAVJUoKuS7OLGXHTxiLMh6n1w6wwM4gwdBdYXAt0jEBtY8yt97OoPso
qRBViPqQhR0InHK+KHRbi2IThDFFRMoiVhOBnBxNhnS3YExx1vXwdYqSoGl8pIQh
TqneC937RHRIOrW7NpnKODcDdFSx75BomBBYhZu5MkquMO/SVLlECgSmh1gB7cbc
9F1j7wbb9ielhfV/wa6k6A5kX53SaFaySY9qfEjqv7d/CWvIGc3+zDvsQkIV7fZQ
sJ3CMAf7qHZqs0AytjNSwSgYDHo+HV/Czc0BODWEoYG/VXzHTsRGKbTHsTxiL2Fy
MXep03FBN3/Ov4sKHM2c89Ex3rxEWvLSFLWTVuk+Xwfc+1gU1uU1jgKJtU3VQ7tY
ltGccPuc0jd+RGse4TovZFUkxyjbjca0bUmc0pNGATeSiEmjNKV11h5rMdgmNdQ1
wFz8TJvKW3FWLm+YjzB0KE0Rlv+4BSGk2807xsPwee9ThdZk4Jhet05pIJMYGus0
fU9HuxRCSH6y8wuzyuRsZarBfkzgdx6tZvWNHZLxuj73Z/a2Gfd+k0fVFj1iR7YE
5cqAUFP9vNGDphDo6wFe9kImzku528AOwJCgqu1jzcRjqMKgfkp34Bv3x8ccJ0Hr
cduiIDZW9AbqeLVLYPLAji9aJBZxhM4T0KSgvjV8CDLVocWHYgnORsaqdS4A1OQF
Q9ghPJihYkC1M7gzp2Z3KxW4ltTRPh6vZm5GUntIkeUmkdVz2xw9g4h7tSD+Rjw9
4RboWPwVwSRAy47YLTwlv9zdMgHQOsOvjlfBvgZb8/1tn+O6kiathyonK8wTg6n4
AnEwjlQPdFrJK3o2UDDd2lkOkmpBkchqKuas+WfdT3eBSF4hxP08DgUYbcppR08A
KnA2XDFBFzvbcD74C+FkZi5Asc8BZuP/Njt9U9Bo8SsUyBlyiI1pIjkrfmSRiV5v
8fzTKFuMOqGKB007gJradvDya+hOBbq9AxEUHfz0Cin/PAD5mEZKxQwXJ7hQc9iF
NB8FVhLiGZGmjIKfPKH3HXohRl/cprrx1SRD51uea4urSkPMOzm76PkHxUKuZdYN
Ul5wtVSbl5h8bxZ10dYiLSx6KC2tLUVc2AgVq6mYiaNUFeXszIal+1dOPOqQPXQ0
Ip7UiwKQdxZrN9elgk3BBs43ynG90HGYdPLAWH/3etQPW8t4OjbYckWeOH+GZZp/
cQGP5op4sVWhO9SbgRO9169/Ra5COO7LfDw6Yy5N/vaAoERJDFFC0uAqS9r49u2A
WG9dw17nfTtRcDBZ76NgoAsoyIV0HLN4nskUBHDWke7dW5P5ktVxWowEpdHtfTwe
FozfKMlNnCcnzZejnkbD2X1rKBVZI1Iavesqrfq/IcBjjBTBP+BOGfCGj37IUlLX
nB8jTnIIaCBq0gWc/vX6atwafjfK2/RGHv6tqb9jrpQaDUjJGuCI/CsIJ1DfHJ7D
llDpyUrQiM+6yk1LZbtloYaT08l3zMUQqsllWG6tn7JYjkcTmj/0fGRqGxOfv7gW
3+7hn1RF9A0L7AjHOqI3vTckcIXtV1eU/lsEuiPzpCU9EgKXgL8ElqDtzZjrEMh0
n02zhSQOkmPTRQ4JFOhzMDRW6iAvenEqZOlBnlwOkCUP72SoDCSwXh9h2EtId+p+
8HmDG0rw1vn2k2vHZTeD9vgl5CyKZjmy8QQ9M0kBqjVuMy/xld8Iw19E7jQWhkkl
clZ0dOP30b1KU4r6yX89MUcNaF/rpn7LVWN5EfkMmP4MckDLBdWVXfFbTXwAHG1n
Ey9cv+XJGQJg6Zj5C46AcpIDCAJu3s8jClPqxfioXC8LCeUsGGHjNeIrZlW95B1w
UWQ5yP8fW3Bzv2wYoKI5eB13xiJR68PcaTd85dIBf1HRxqtkgJVjHzSibpGrsjgV
BObyVpQG+Uhc0Kigy0pzn7nWQQVCyyvAJeMHbNTNz723lfWDAbi30t4QNpO3goa+
e+o71fr7drbYSo+4SFQUdx6+sOKQarrN8YhDk6W34laU0CMhfIgcC/q3QRwTiSlG
nUDy8z6lMBJ2bzib1pq5lz3iv1suePQEaqWamFtf3SwPBsLPryXtgfaOyAKBJPlk
tJjghhZ5d3YbFpB6ORhTJcg/jE4ol57Pj+r+GusE6lVHnwXt4C/5XoQntYcRzeJu
LQOqN6QjHTEly2WNm+e0HFRNXj/h2PJd94EID+c++yG2eosZcXd5oICZx0vgLKGE
YgGJla1IV4ykK2qLhfy4h6hQzJ2CzAdb3jRdcdHs/ePCkk9LuZIjjiTeFxgUUssh
bFtmlcict5QoobQwnED2tmtkh1IV/ZklzkQ2MvEQrzz6TLXEv7c6uwO4rLcZ6fvl
tjKWtrVqBc2xeNovFML7YpuqS7b8wKyRIIZ0XT+YGXD7hyGufNz+EdANou0R7lnS
A4BmbXlbSCNVHFsVb/512XNN89p0Z0Hq+rRy4pue2X9sYNpYMv6VNm/B5iJUhVWr
UuKfSKi/ibUVxrQ3+9kreX7/Bq2yEmaovhiwKBRsGVdsJTGHDf3onga7VS1gHnMQ
39S0O8f2Haaoouy9AxQ7cQ7KhTLO3JCJRNxbQEh0/ZZIHgHmBB16QqoBm/3Vz7x1
MIq5b/DZMDCNAK+87vTx0Ah6il/gwvZMNkecRpBG5wMX9g+gF6ZM1O875QYvpuwG
qELpR/YQhKaLVwL5RekIYh2QLZRk6IP8N7EmLBs7ofvePUlVRIpJlLj0ab8WwOf4
sdtAADxhk10TifHU+1L4kZlqN0WDeJ113/Fb8UhQgM96HV2qVVxBX9671u7VVl1U
knRrfy8mHm85Rvoc9C77wrfz0IZk2KcbPxA42jYe7+EggCEjLVMZWU04+Sebalms
WXy6wvROHb3Fssf6kV4z+6MW5lBJfzJEHoXa4AMHcsY1NyOlMbh3qJe8VdeAHrMH
4ZSV02KDr3+zc5Rydr+KwIF34dBxgrYdwAp68ayMDVg4gRvRLlrZZUVE6uJhDAVw
0Sre3CfFp0QTkMd3fws10MHX2vcAyN9PpQDZZzmxwMbuiiCu8c6XbVjT1KwH0yap
brQCt1rXS8xwpHY429LUVZd+QQQ12My9x3cp6mipzclFONNqtVeFC2fw0UGjGgmy
vqk7VMq4LFzCMaBZc8MIpbIjb7B4nv6RQiPWmSmVSAjftBy2Tw5m4e7snpQeS8uJ
XDUb//3EPlq1gETyyklYvuhfb423otFLzhbYXhm6nLOK+f5jskowYSxKVPTM+uZP
9aKbyAcxJbKrq8Zp0IBdsuUj5NqB5KKTNv/9qHTKj96j+vsg9ixBVOWAUNho8S3A
pbZHHn4+CePbBwpOmKvCeaFveZmN51mQyGwKU0XiaEFbIVMNaw05NdaAguzR62At
JjNj8Uizw+q6ThYa4UWMX4hV7Rf9GC8RgFeAGjCZWbKrRyvw06f858lUVcSq3xLa
RNO01Z9/zE/3nHS43Wu4aNY6ihptTVCg1mATPMl4lD1xYz9bw5Ze253KJVKrE2vC
DVAFcQu1eO8ej4hoIKPy7CxFRu/hwpaLLYf9FcBTKxFmHKCjHgOz37cWHGwSC2O1
YMyMoKtlEFhGMdv1VPw89UVsiAflYaKb1V8Kn4Y7nYTl/lchsPXlh/Lh26i3Qx12
M9dxF/elxaDGOpdbVy8sZl57izpz2t7C3ScMALig3O27yzzmL3oIquJglB4ek42H
7navmWwOwDTX1Zv4Lfbmab/LbyL6hfX/LdFV3q3FsnsbswCc+KBs5zKMaz4IWQ2x
prO+zV5P5cucvy3ipdiBP6AlhvVoXdtOdCF2RmKy7ollIrH3NKpJiFQStdywgzNR
zC8mHsGtKiyFpl/PEkP06NrWac6v6h4S+E2Wm7zCPipVAsf2EmSODX8teeTZs8uP
wS4WNUJV3QaGpC+OyydPBhBmG3mmMYoA+/e0A9NTfWXc5ahUOPckeIBYi9FZTUMp
CHiqnd7Fh6FUDubSDbbE6i+rg6wlk6Eee4PHNawlX5Yz4uy8nEy4Jh/xn2GdWtZf
qHBjnDSqxEdAujcBdF/WvsGJVZPMvlIjhFbvVzODbmM1Cjh/SPxnIuue/kyZRG59
KID3CJCaGWvSeBhykKzj7sXj96CKnQK5DbA8pkzmsVt09UitkBRnbUCwKyDbEfTR
S15/dvLSnBOdCohNSLrl2sDzRgBTATKlLtHLrxduiJk3gA6LYdVh6zMWVge0vdFX
KWIY0maOwF/Gx0oJ/rQzpU+KsDUGJths89ZwNQmY+WZWDc5K4m81xzIChAxhu+0p
bgDvLAR0rqiV60oZsX6msaQ7EIoouhGGLzeg7FDk7swczGl9a7ZbLF3020J6szho
5QMsiAR/k7KhRAlst7UB9/zQ5p3iaqomxO0X8pGx5eevkthaHUqrjlnFcRWQAfyf
vk8qSoCn0FhTaE9DO3n/c5ivnPrARuOUzP4zROLLAK7MCmUHc0C60FRBUgATjjAh
GK3LcC2ksNs4vxmvqbrpQT1F//cjA48pQRk6KB7Xv8J1QUWPQCOctDhkbX5spVTK
9ymjuYEXD8NiMN4aNnH7H2BcB1O7fh85auVfQC167jP35NPL/6B3r2XxYlblCd71
2rCPAguYNS88jUpEvklUZK8WHAe6nMNvVCgZJRB0MLXccPIdC3KG8G2mvmk3Q2Fo
f6arHqHun7ewa7LH8Rll2Heq1PioEepo2kJkbfCMjtKINB6VRMtPZxx4UoTePLSf
64Kil8+wjEf6aqZZPLSYZMEjlp8/qvdqT7tTnDgFU3VXsyFM+aVAHlQqmtwChrJf
Dst86wXm/t1yfTS1hsYKuWOvdfEWceSmJqajCGuzIEhtfigXCnuark8OsCrwngn0
V9sOcttlgbO0IU6FyVMQQykG1TTZGaBqoxPxGVsrW3VNaSor3y3Lxkscj4W5uK8f
T046D8spyvxaKYqKrDRTdmGou445Bq7ETsGInb07+e4WpYF+39ZyqULjOGGHJ6wR
mdTb79pqtcXlByVaBV3HOhEOxqeiEOVH8fK4dgxRauSHXnaP/NHBfSG1/21P1q78
5r4euNmqvQQjiHYkv1/5W1d9eG0FzMBE8BsxxLdIOtbkWTb335Aqa5VNIdLMbSz4
AsqTYCJkUWNDHEg0urQGRiaGe+H5/sREHX42rcP6gKA9xCjlfgpnNEW04czKR/P3
T6MSXKBogAffUkTxMkfSO5OBIUkklYlvpNquvjt8pAXVBNJYVdKJhrCJ85dYq8Qv
rsiIo2QRWTmLo8Bi2Et0Anaw+DO2ZcDU1bhotrVW8KgbsmHDizAJ51XfiLcnwuIo
3LEVILtMsG1gGVKIEWDTXLNaPAp0KaXg9iLlHB+BuCZ7PSr6aWhuvomg7ni0/eML
k16dNo5WvLdpSBYMq54yEoGbcaDFcPxt7svxSn5OPNp7xgYPOtTNeyMcPy7TAA7G
cblyBTJpjXOgjAc71/nazdKDFSXxu0R7+6S7iusTdcFPTzSAz5/MrhLm8MDkViG4
24eFaDsGblJ5PXsrq50f562uNVzsg3/Knofq9xnqv+RPP9Jt6KZZpKn8o7/Bew4G
DsB4SYEzc0G6TeYRoz/hScYsPUyR7bf5m3gJXupFQCcjkHnHmr+sX4g0PijSkFnW
VYjZuSpP5jUiPaCtuLOZ1IV90G6JSPVakqOtJVcTxBfIs5lVT208ajOpVvVQFpUP
texVqPZQ+PM5TgQVgiPg4qoUmrYEy/y7vuLXW5r6IY6gCFbLAtfyviV24vawzeta
mus4qW2QGoMIIG75earXLdzVMnBkSmkGa8oMdb29y+dG77rumDLKUaSz34VAysaq
GMSl6FmA9EscRtCxxPY9U1esux9Ew7O6cfdGcn5CJOpxcgtG+GDFhQXrvcxibbz0
bPILaCeq0hSlTMf8CJmgxYCbzhk2hJadE/xDBzFgvPHUeneWSthPYqoCke5TqTLC
e2GQov+R5cjAvNvsFyW1JRLXiv1EVZ+6QqHwMWoVbVA199bnWxDGX0C56kZy5AEv
OzDLEzWaH5axefncbI7IZ3Qdua61cFsGf68J3LpRbiYQN6UpMOQ8b0AZlNFx8rRP
h2oAtqdY2xWE/9zYkomz/uRk0/u4OsalVV/Dckh39ZqWxEj/fhFcmENIjyw/iIof
nIkOj6Gkmowqre6qCYyTUSx8OCcJeyJiDrV5fL7byJ25mDQdBsc+yocQHXi+GLCJ
rAz7rejvwHpwY0JyeV7PNGGpl/Qw8yGHiizpl95DjG7PI7psj0ZiGuz/DA2rxfVU
epZ1mD6/AHsRAMtanOPasoU2LUawMe/lTjcvipzFb2BRH0JUFL12udwhA3K8EkiP
lshOvg7Eo/14Jk8R5ZaA2kvi3jElCaxwTYtg8DOyE2ejmHYJAwmff5lMjwy/fEDs
e9E24i7Amb+y6GW7Mncda0FViXpYvZdhBbIUI9YaqdK7p8D+6GtzXmjD5CF6RT+7
I1fsquESrrRTxxkqwzMH5aKq1zjQkG+FFk9HkC4M3vN990Abo5SkNi4EHClspxvw
HlOVySsXjI+7nSiIkfq6E1jNnQMV+EU258MSohyqUolkSLSsMnUmn1CUkkzVVu+g
gED2XmIU73nBle75z++50TmhSPHM58InmfCRzG2G2qU8WKDPL388cIzkCKnVj2bh
q/A0lYQgSLm0dLqYYrneA007kf8frMX76Wd0njCSfufrWdFCOOmaJWbQGzNHTjM2
CMsBEtosOTZbaLgJRtx8Tn0kQvgktPkFbUbRgZynL/r9BMxn1EwQTRagTT0xrM8B
yzzAOkXn11n/mxuMBP8fmQo1sony0+EfifiypQjzpmQ9DLJ6CAkj5MbytlgZxiwN
9mglAHhSqyTaP8h3kwI0GQCmeKC0jMsnv3g22Codr2M7zOAnR2ofkaq+yUBF0KkJ
z443doiKNo40PKIF+isouzlfwqo/ntmPaNc8WthW0i8aIOaNXKmaemmx2BjgHBdP
l9T3TVH1My9QO1VyYXJy2xb5IntCN+U996V7KMz2pSWz2n2Udf375lqafgOAZFNb
Pe9RX2l+EEMfpTL7i/CxTV/UY4H5pMHP2nT75ZFxenTf2rLz76znoVud2OPTBM+4
0m8j2CSNGXmSquLGsG5BxFzCFH8o2uwY3D9S2dZ6xPHJM45G0Zz2PRXlsAvOvgvE
RpC8LzF7Cf1DxuKI+05ffyB56gz8sEC+2JPh4zvzR0ZBCJ825KNAnCPx5jEpa6/m
PAuxuCEqQgZzBUJpCnFDKxc4oBIr8N41dDfFBbxl4DqrzqrD/ijuRykMAF8yzX1l
xFlDf2AKR+6mGktD8VEALeTSzU+ykbuoq7T3zeLDWPQf+z7zGyZgrYmu2II03QO4
LpH0w0Kw66wv9nrCQBsekPSVexgs0W63xHOWiub6jOfpvB+ut2Tn+D63PZ8BvoIC
WZMoHJTUzWhWFmdWqE2B4Y07OxJlH4rTu8/69Q5DUvmEGXeOn3bCVBmYKGZavC6n
i9/Vr88cUf8G4JlCEKM290ueJyyzxD/2FaBtmPaB/a5wlb/hd4gtOaY87LtsgZrW
OdQMSHUa298u1PrGG0kDY4Dzssz1MoQlFwAG8v8bz8VbUKPJmUy/9mgy81p8awqw
jf5GNEm6nj04tq463nyWYBOAp88BDKpS6mg9WjUP+q9MHqe42X9acpVhqMWFk/5W
yFKm1wc2uSovGFj0+eh951vmKYR2K9iP3Sn5rtHwAp4dEMyV77ZJS5QuZFT1ChGL
+O/oUNoQ9ssJxGeUujUqsU8ivSe+dl4juDriKpKUzTfOvSUl3BK/6H5lv5LRGrOp
ad/4sqCJNQwMQjY9at6b7Osg9u5CUcZkMu2HosASt8zXyAI4i2uksxOVwZ6DsxW6
eRCCihN0Dt0e3CvQI2f4J5aVrg94UuzpTztUnJsT6uOneqL/m4fQn59H4kk6Tsjz
DmjAF1k+/vAEZFrEUlg/Nbq7dardNLwvHAlEVAGOvPgD8p/0Jt//j5SdB2aia6FQ
DyolxVgZ83v7tSiRE5aShJw6GKhx5f5vXhx+eQZ47tz1Nt5gmzhY8eNLUBiVWF0N
u4weRtaUZHM1GUo1JLTL98ka5Gplw4E2Ce/LLJ6mzUoXv1EjZuqx0HoG1Ug0Ky5T
Yz2cB9O9C2MHWZhlZb7BKPrEHPUGNN8mKv84XNhe1zd59qMcAWH6WNfuK3eOgWV8
gUEUZLkwI6+UUNUp9Pt5OZZ5WqPLo/92I44R4d4okOmylccDua2jzHPNtAINb42H
TtleMS1M3vFHLislTvhCgM02p36phzL5xHbeIO+Dhl9Awl5ppT2SmDv+EG8UrTfY
0UfUPhh9c1Pu/cG9VDzuD2v2ukreow9h57AmF4zCuQEUGaIUbo6x6ggeiEQlz+XP
t6mddwGGCfgT7tySRiFhBCBeZISXSRF9DpO7evLCUOGQvdFpEyQNgPV3JaDtBmEA
ulHZQtb1CS+/vbFZsIIcLDGvThFeUdncWRznCXG7F/LsbFgZVHbHZXnFU4ATIFdT
lyTUjPssd7y5isyxpLd22PIEfbKisdTi8XYpgFmM/E+oEPjmVNV2rKZsqrbDoBd1
ceG4LbOvm27nr5oyKGcvswDY4makT3FO1bY+bUfxFyeSq+CK9DpN9Odqi62M5GOp
igaZOczs7uEJTcn098ss0BgArXzSOqatvD7hFiXTaJWA+1zanywLy545FLa2WSs/
u5PWhjhKYZr7gFSziMB0U6NkiDFAX4xgnXg/arsGtLaBHFWJJUavUa72Xv8AkI3n
WZ/uOML1SDEHfbDHaU2xlEi8aPMjtM1Tgn0DoqUQlfFDLSLH22uEev0LK95ktsjU
xGKreQXLn8sg2XI4joMu54PfQoGV7rK4MoXC5VaHVEMaWj706JZJwcpCAUq5yLCE
AXL0NvPMtAqcRmIeNk/YAvITLsozBYj41MXhAvXLNUm9p8nRZl6v5Pe1n7zcPsUh
XSalNbXiGqGafV8lfSGfs57kxswK/YJ6Vu91/IH1IrD8S+DdkuQ0tf8hjLA2iWUa
abZUXhjTV3wRBh2qdpcVe+Ztj6Bm3vjWU7b3xfRHqiVh4yXvDNG2sbZiLlJ7fbF/
Fe6uy3lGLSgwZAWke31OgW4aMHPhf2Gia+PiahQN1HZvBDLOtFQInJKK/uK42Y7k
kzWsv5gB7xsGfN8iAYM/5fJGUDUnX9YitSOS/w6JHpr3iNgbxF9qVF6pRx6O1vTI
UVPrOmyB4dYBqCn6+fLYVaRi4Yb0anFyw2S93LAIia25Kp85MGJH+T3KBYeKThPK
1WZTgsDGrytdP3aPhlv124KuK6SGTf8QxiNet4q38TFzGwuUdrxKXkTlgT9CdSp/
BUzj2Rchw9L18wOVrvcmaYd4mT2v6o+eozMnW4HfjH2HTUXMJ0OyeJr5aNQ03tSr
Q95+sISXypdwmofkO36rxNnUnZelmQB1t9zNfr2ewcS8Ur/pUAjirAqq5DxsutQ+
Q9Yai5G0or9AM/wEJMES6jYJrghcAW1lnIGENdHZLDA65wxktBMIpIkrA7Mvz4CP
LDt3Eliw6sp797itXtUrfpFTGZSjGx0iygSCjPP7TySHOrXdSDQimhMjvbSOkN64
FwVa4ZAAwR5X/p69fnKH02AEUbgpSXKSvUsTmTR2N7f3LbOv2fPPyxe06Hbu70Xj
EE8Xbpa13U4qFFCoa9+Yr4V/WiwvF+fs4hOJ5zv+XK39q/sp/cWvY/Cqa2eOycld
rkxagWoFBN7FP1XD085OU6ZgmiIsLGOqRLFyMoc/9rThXqLxLWtinWS5gjmyoSac
mAYU5WyS38fcpztG56S6PjxkEyKXGk5tK4w/YB32OQyIMzXjyuc5PmRH16ffZiME
DLc0wmzc+D5Yz4d0ZccWYB0hxHpHEaRTF9EMpd5MdNGFwpYYpFgBu7O8M/D5ao1W
Dn9V9grmK/s/YbqGi3VfF1G10T+8zJUHx6f8vo5W4iEd1/Dkx617WV1lPVdg6rgf
UXsx274Nu8bsf9ERyGX4IcGVHgjTag2IoeJTsXWu3fno6kftx657RQSZ8yHmJBqy
9Qsb8qODjcS+HxdF0+q2e8kOsip2Sbz0AxNL3DyYzw4cbPKb3ntnReGK2PHLMLlf
O6LKpLa82yUOKIPEm64mmnhtLWd9nmDLO1Q4Wo2+ugOo+xW+Aw2T0guvs6zGmd8Z
aryl5y7UUJfSF9Zp0+YZWnxRQPYR6ELzOOmkSDtBbdzPsuziZ+G2YtAk3O1A8/Cx
nFA33WRhB36/u4fjDM316NvlixA9Pf7J2mPEtZsmQ2p/l9pUb18rw2tWKdjJr61A
V9LRcZ9p4O4sjnVTmHC9XH2SIKXP585PT7dge4XD+0J/xfhmk1Sq4iEXaE9Mw/J1
trOBarzEyTDSsL01Jco4M+5JqAU0XW8FxH5nLKBMZzRAIrw6YAbW/u3Yt/GP5iuE
zVpemU9HUPB05B/9pZeTW6WF8Bu5WeUSA3BDwEKZnn94087u9SuoLQZyZQp91eh/
MjFLSZ4iyAOHYaHX2t+90iV0Tz5M0tSaJSIQy994VvHfy5kbnx/zHr/dGl5LpqdN
3yW1YvJ0ubjUA7hyZs0EtbVsfpWdJudDzBcjV3+uOVw89kTQKF3mKRfcqKiW3qbn
ApZ/4waV6O+s9+Hc9yzFv2+5G2SOutNOAPkJdg0h22h0rHs3qDuDXgfeWpan0vzd
RYNYr+CEu8bqYc3wJdLIa/srGCn2MYxcNBvLV0z2UwXZ9G1K09LiUHNEWJh7dHYo
7qW4XvV6PaDbRgCdhSvazRNKSHjiddK5hHR15IsR1Gtyo4wVfCgwT+2pvzoqffjE
GBzH6V1b3tm4ZFhdMPQ+hihzhJyQeCcp4WkjcSU7wHxtE1CPuY4CCvFyuFLE/+av
qzDKNOPxFqddaYrKiPGkm8uedYZqS5Xb3+rf9AqfB0f1X4MfwWpsoeeCfkbnBaIz
CNToxBn4sYWrnDS1sjzn8HUOpq+5BQlrUpuDPrfmGDrKeXH6ARoEX5XJMlAjMj8J
yYMjOus3Lrwh9u7JlYJZ4AMQsRnqtCdQy247MOppMM0St9ps7gsJP84QUhMMKhAm
TBlZRIOPgcfS9HA8DanecFGa/yf+Xk1uBsrHWWwoaZfUeEftl6vpdD2D6yzX3fAk
itN7rqRMcQslbuklQKI47dXYf9Vwel/IpWf9ncRw+4BV7d1Q2eiYwr3pGDelYENz
vK91E6otSDzwKbIkXdxc8vxD6D6FSZmQHF0b/UGvv9FB6Nx4t+O9UUYGFtgch8Za
RfSS/3qbIaupR9xlMA8c1mdvUTBqHM7xc3oP+LPM/jOLCSoDDvH09sh24MeCZ56R
+PDubNZZ+FOUbqDASWxJUIMt0JjQM3P+2cNtiO26wKOQJRbN8TGqQKvXEiT+uUEf
4rzGwEBPpTRu5C35IQ8H03hb3kRraMcPIBdJUcpUNM+kBIzYGn9F0jPcSx8oRp1O
iqXkfl1uce4Sy/hVQdW4wpOactf5ZjZ6w6vSaGbgBphMVcV/WdwPkgzScmYqQ1+r
EdXWuv8w0NELqGqtuHxj42ke5XeV4PxEd8RDMWcLfNv1YEJGSSPn8wO/jLFclhFo
AGg7RLB+8UIqz1utaIZQXQlA7vNUYZnjOjaXzgy4gJ3uOwXvwfImCx7F3ZI3oB9V
zoKZkQDmnHgD4VztmSVLX/a2G84d+45sznt6UgoQDsVdZGAMJYd3Q7CSrbMAtENo
SqP+FBa1SggiZm1AYZfIAQ5SM+H3+U113dRtUhLZa95TEEx6yBmnR9hruKwnTARh
AtDknnKDL65u29yGGmilCru0NXGsZdgoJ3iOpcnbXYH8mRf1gW5tDs3O1eZBjZV5
pHfXRSfJ/hbigJ9gy3iHYweyqgbjAT+a0giv5Ui7DiCw/kJWk5ih+qohTnjhsskr
Pt2gzkLPLdxX8MAgthgv4L6WBXC9pOgLJeLgouhiF6C7BquLV1ZjnQzuPe24khUJ
UqXCN3ZJTU6A38ndX86MZoQrc7qVNxkurWCEg3VerFxlMAz0oj3ZJGMuYV5fn9/Y
F/JCv/5OzvNG4QdBXrlwgZjATVMGK3mkqDBaLl45YfSj4FNrUrT8X9zjd2pXL8bM
vXjKHApa8WykKDEBS0j+DsCZ1yFUA9b+pxyJE8dHJfezky5fUk8gkKLVLEK5jFNt
xYMqqHxHhCP+YOTLs6Vcno+7T4wPLfEtGruyZFafWZPBgXzuhbBy9ZX7kQTdq6e9
Gnp7YpXvZLyAG0NfapE6+npmWT+jo20LjlbvK94UtD1YGsK13BIj5nd40GHK9AuU
n+Z5+lL9+me7PYjXeVeOLo+DKodIFithZUCY8bHXVKzjVPb4Cp2OEjnMzcmbcJIo
wKV3JzklAxc7BKRQpSlJ4yMW+K1yMZFxPVbAGgjTii3grTWVLSryalBEOXLmUDAG
TQnAFfv8XpYw6MNd0TG4Jvl312iXuMUTTvtYNkfLlpE2gL/rCXq+lIWFf0xEmw/c
uDZidlzWtptLSTFRHKKaK2EcvmhSxu1011e/sYW5zR1mx+CGT1U0r9AW6Tco3cPl
MwzD5DP8ATRwB1wc6x+n0Q3Li8jkOODk3MRuR85el31NsgrrjxQgkKSGBNHa47Uq
8/McAe8IPf1HOYwris9/eKCi9v0Eu+qyO2kABxhiEtkBM6IfkN8zi22JBbMUZYlq
2CPWGpXfJLHER6pysp4mmbwGYwRgfV4d55HTbICwE9hWqMSJuea9BLQIPai40xch
iKTUiq8Y92kMBCY8EpFKjX9gI44z4EOZCTtY0mK9JI6msHtInKKvD/SbropqB7Xw
mufNIFgNG63eBy0PJxPmoImULHa87BK7jL1nmHUjpmKtqaz0wKCakvPWczFwgspp
ZBvyAdl7zgHA/k5xoepBl2QC4SdAd2A+UTQZS4Co0zYuPLoDkqx7RgsqUw7/T1+4
f9uTFOP+HqR3Y/W19W18qRjFeexA65xmYAc3BRxrsP89NjMFIueKhCRiBETn4RoM
LtiNFAIelEC9faAxBJfPGG7herJZw9NzXzteg9u/PbWX6Qz/c9vxvEj9e/APrv6Y
EuBuleEKEtCC9pE9R9S/nQwYvbtc71f4jv0N+hC1corj5KmVlan5MIPArz0u9wG9
BkUAnC8bq3w99BsqXUSSLbQNhFFAJcaUS5EAq67imVjxTPpJxNpkWuOqxFSelm/4
wRsaUZvS5NYr4wvxPgd0Qg9fcql8BfgjrrNTYcqDBs+FnH5iQFCyOo5TRsVxFDBT
teDlaz0ZP5aXB1smYi53hSUEmt22fGiWALhLp51dGH91v7UHKmLHT3HKZRTjbP2R
SW1ilJ8acBTMpmjywepjLBcqkWwnlffrAN+oOUmd/DfHvJnoSv0HwOTeHoixpBcz
9uKKXMTTjZaghE417Eyff1oWrouemKipc/pdzykE4nqgWaz+zek3lvGuS1umkxI+
64USEyByGwou4mztnoOHrC+ieFKQfBCivSYQ8W4vvC/PC0d4+zpwTIigwNGQOP1t
d3uAzvjTVtPCpCmd5LKQd7zhdP3iDiDIrg1EYDNy4s7IZvE4dvC801j/PhxcS15K
CjpmrxN/6ppMDQFPCgy9837HL0xpcMc7Fy3x4/VMkPegQQwotHLvJUb16KS/fsRv
Mp1cUPOCIUZKPY0vM2NYk68423hA76qvz7Uko44hBdFKQo/bzPVy28VGaHfGyS4Z
DFwYPipavW9uDrxC22gb7sJQzKtSU/+uep72cdT4GzhNCW3PjbYCPLl/E7bxuYAX
3xxbwelAjVy/hB3cHdhbzYNY8u6Tw6CM87p7mxJvYtnSiu0V8PcmCU5Lg7A+IAHe
IwiyAqJHZLblewqWIl7V0Rdus9dj9IfdK4B5ntoj58AjQ/YRID3tF7XwxS9L7ifA
BeGqgHxa+CAeSD/ti6ChSWfT3FIwm4BTaE/75zE/tRZvy14Zq9LmybOwS+gtyFp7
RSawZXZ1zRQCzlrzmGy3OjdEWafrOn3e0oMDBzi2lne4A67K/syD04nItruL9Jyb
O920NRPF45YRGwgqwK+SJSvOgI5fBR063cY4s9DePSJrdYzUkEKAd/H2G056jmkf
xDr9iOJRVPsQOnrc8XHwX6OB6xRpxUiwvcn/BAa//ldZ+UmPg2HBOFSiGXIOcZyU
kKbnkeLN/gozQaovUrmeWrWZWlU0+J4iWKSVnIJzCbZh63WYnc6K48ndHVjcC03B
oPua8o+pRXLztSgORxQJAOauCuSItC3gqkSl4z0wrqQXWgbLCnkaXH0mkdr3Yht7
M9n38OzrhCQs2UMRLOYkxnXKA/avl7so+EMfCdF0Ye3Y9JETVH3kKrbZeJIBynQp
OVvDeLOvx23WtXt1NbHamZhEJ7HAEV7UiPYcpgESlS6fny3ZdheO8o2aRUuebK3K
At8tPhLC1+em7KVaW1FDiPYupVXOLagLu82Qsv6mBbiteZpRW6SHgABMpx653F0e
egMjx9dCqmBm47HnrWp23FOv15Ex7TMIUsfyAHqU/nR7f1JHfAlrD5RddYUawF06
w7Yf7K3zdhJVB949B5PBijrEcn76dFP+EXzqbGP97LEOVZ4KYccJAXSBGiAscAnh
uZ7XhhEcMuqfMbY1fNznAkewZKeLHRS6y6YyxB903+ZEnr9GUpGAnX5tpd5XIllW
0r4Ejwt9BE0x2h7B+qZxf2dBVv8NDXvr4aModIRN06qFcZqW0K+1IrG6juzUomeF
MkhS1zdqudRuSKYZP/NETru9FP2jd/wR+c227TSO1ZDMWOCqUd9RaIkAv+LObLaC
xhgFwRrcqLcyoChYIvxPcn+FBuSR2gbq8FucbqPEZpzdUJKDX24gJjWNDx9JlSBi
jNUynMs6ERrK1PKbqBX4Mrvj48t8SltKOsmskUDDbyoA9PGaR8PvT8Y1QC+kMdsl
tv8lAEXWQqdObq+LvLQlX13LVtqaFCVdx696RISq8Lsk3Omy9p74kfg3TjTeVVvw
45TA8VD5SDwnYkjNGQbilPVqzLKNn3bddxLIJ7xKGab2PvfHhtiYiVPXeUnsCiNY
tBtTFZD4+ORhVoRxhYD8lwXdB7YmW9gzVFhwPFEQyor07qAciLiTmvGbJiz3MWZM
g6RFzLduEUhjvENqfEChquziJ/DQKm/x/8/8kpcZkDRYIx1fUv7Ztp+Hz+uI1LwU
3CBphTp5VFV00j5k+UpWPCK4M64yoP5o32cBCxBpgEkJk1w79hLMFhCneW3/jKg8
VsC8ai2v3XuBVJQxP9yi4ObT0/4QmA1GOIHzYPj/G2sVzcWgMfVQA+hZ7LSWKp48
KoYC4uxA4JIYCwnlNJESa6uTE6vVS0cfDqPkumRAGk2+otLNpV4ItfNWpB7sXIrd
dtwdi+Zm/sVZvRoUSc1Mm1e4XJRoiAuaCG7XGwUENe/TpSZEO9M2DgFhokYjyHbh
orOUV7SMgIHXdJWidKbF7c+vRq8O05NJ9HNMcicixvPlillispJAAyAqVkElTvdP
6+ChLBlMSI/8UCFIOi2YxQ4mlfvRMAp/mehGzK7OkIY2abLYRSnMMY3iRKnzZ8dP
N7UMievA3SdMUKS9lwrjHOqWEjkLV64EAOGpPROVHpAQWw3f4gU9OzXlD+6zUcXR
pLig7cEVSCaTOXYhKpjbSe4cV4ThJCBJUAhBQ12mlgKzZeKPQJYBXts4QKgxFoiw
NalPSsw8TP5R8CG4j2eQT58wz5LElapv+jDEcInckY48SxdtzdmUZdvg/PjDpimp
Eun0iDrqYixCO/228AWgS1Xa94bUTsK7pnEqX6Na/bAjiEXMUDa4r/ZY/xgosk6i
BhBjEILGT2S5VBjy8O6Tr6Ybwv3AfGas2jkH3am89imViVDdNDPDEIVDE55TXJ9e
FnHx4FTQVE0D/vZcbPaTV0wKDLSmwbYB/mQrvMTG7jxIVbSvQCoBzitx+DATuaTJ
BtNA1D084fe53uyd4amCpBe8vKHkky8LZP+Emg1thLApulNe8l60IJ4PstkgUb8q
7hv+mzmIY++sjm+ENNGcY1j9Px0Kh9dhEAea6q3y5BqBcE6PFzsFpgE6Y4Jl4rnT
HP8rqd5KfyllCNkXHU2SGpImUkicC5MpXU6dC0GzdRirUzCJDZp+7ZOH8kqPLeXl
i8bNU4CJu5cfyMXdxy1Ni7wAonwvEvKt4ePB0KObNjZTm6ZzIrxV1anMZ3KOjtef
+RClWMpZLF3VPke4JLvNMfJ0+RTCmNMJXrlachaBpBIZ2pjRIPc83cldB68vELXg
w8tMbluMco51m6+bO8R8SqwG9oNFzP++sIY/iMYkcn+juVd+dGeMiSUCAkm58T3q
QOF4HznpuTeBof8oHyD+cBZ1nhVO3S+dhErj4XctDftTy4TOQfHsOiKhENxE0LBb
CCoJaJYQcAMvrxjcFuz1FMAawMqN19cqV/g8hjrClxxFQuvRWPXogoMc/QbIEv0y
7ZQP+CrXKIDU01RGcPHZamyWadkz5evV9F+0iFK70/sjy9S17t80FsIVMHT39Vbe
5Xc6A/bcdU8yJyWNDx0z+vV0U9mczesf4uhSLTi9aLoJsFN53M/CO6edOPPB5BZm
tiUyc0PiCZLfoEV2XsgSHvr09GvCAUcGtOhUgw+/nAwOfzNday+cYlSe2IrRE0q8
6H400Lt8jnX3cowHTNF0pRVf6W7WKxnd42TbHk92mYClRryJ8/mYBgqTOXe8hb5D
UN35B6oN7FSys04xLCJZKEB54MRIN7DWXqfRMrXEqlzNazVBSE2ij+O9wPd8ISyi
h/BJOFQ6xumvn9iR8sLF7CVSdvycyTexTYZUVtT6p7zBbbJH4j327eI5Ue0vM85Z
0jcZfi45BnQ93j4XYQlkvF8xhWf6igEUCv4YuFF/XnMAiGwesWo/GKVKHwjhmzoI
l7zFOsJYw5Ld3fIfHou1vcyY/hZ/BC105HMQMJ5HDwooMQzTZc4DrcAIp/43I9aj
dOTaLTmKkkLhCVZjF4FoNoYikuBZEUsUye7BJAabFLSLpgsZRAF4FGsMRNa9kTHr
pXjmuHIDUwEZOTcqSvIQalWWqEsymODIObssNU6bIIGukGMopz4eLBaH866eILOC
3LomLwEiZgoI9rP2NUQ6cxwJ77/zMN+x6HY1LgtcRLzi12zFA3iwzg/54Y1rptds
ED5N5JX1gE0rBRBx5SYLhoovYlWfynl/Nf8703RneJNtc6cAYvRweWxdIqx/cENQ
IYYjQFckbqwt80EeD5LVDYA0XfdThJoX20LrbJZ2CLrtilmRp9LJapDK0L9eqo9d
fN3ZPsTy0hkNgKOtB3sMUu5M6hN+V5tCs1RtOqp4JU0SlzuBagmxnw2i0lKbiB4T
zvF/HZULQPdDkt8L8ah9TavkS33RssfwUe+xVPGnstJ0IhwFj2jppc9Lp+3LXIjx
lr4mqcLJ9VVAebuSXN98CCsNrBGRFfsAFGUtTQvK1wXOMYrW8qYrzAeB3KU8NaV/
vz8YwksTkKkAQFLpeF0Ef/h/Xg3sKuORHjVU02ZwJkbDiBzcUWq67sHuhBtwZeZq
gxHeasJDcVJefGnHkduE5CbZD6YsBIW8NKgriEdNSEUBfnMmkItUTapNPrFcI8om
8T5lzaM0pZpGX30tsDnihX8XtN6eRCF4EWFwoFnTPWqoKC520vUIflep1bqS1I8A
2uZUVP2FmrKYRHHj7nnPI3697OnLz28noeBFlXW6C7qFwBPuRRkRQ20IJk7Umcvo
tq5ngUqmZyxWBz/a+2OkG4Vfu2Xuszfjo4iTFNlajvBUofyyeWPJKV20RYJv6GA4
qTzNubP3IwWLyfJF1yDJXldjv8JnS2IdMMYWiyVsb51RujEajiGP4HDGl/78nQ+j
emUEWQB0HnRqK4O9lrK2Ks1zTrnLSNijKq4NQPXz3d9jDGT0C0xIG16DABUiyjh+
SbpiXK4XAztf78Wfnr8DLwlDo2a/DR86xDpB3YuLsbN9dKyPBfVv8vZfnlXFAKq5
HhGEIN2q3FxDDcrVUhCF1wKdmpvYbaRNAcPqT/ePNpwGPScuicrENxq9/vJkd0IO
BD2G0ZEcK+d8Y4rZ/N2eCjshrlCzI7HF/IAsVWb6XJ82DuaoZvUT1UpEP2GwYnvw
RCN27cry+4t/qelt1mU4YxmFJB0uIbanJ3buM4q2CzsJ2zmj/xmq6H5pBWUAY1tB
m+1l2zOjOuqhvsnwTv3oJOQu1TOvGv++ByHYhZmrRyFrb24WTnWcidXSFW7lmQxb
QGdrzAimDOh51aystyDXLsCVoW18m8WUdEWNSPt0deZf6g5a9m0QjsxhjhSPXLp8
h244OmespqpQaG89nic9BJYL7nim1Fxd8RhJZtQMMllvrniyeR5rhO/gOsaJEVQs
PysUMfyqqp8/pJgtthNs+uNIA6mRRAm2Ym8teujb/3kzby9kdXvw3fuo+SSt5XCy
x5h0vmB51QXhBzGYm0HNWwmud16E7Tkwdseef9G3bM5y7mzzyBSQWSk+4TFGQUpD
3NNDRVyX5yE9of415b6f+nlkPknvTSZKPPm8K+7n1e1gCNsae6/boX/zIDU3KGfC
58olpUHW3os5NtgHtVogjTUNHoYkR6f1l9LHlvBorqF2CfWhPOm69LGZQmvXiATL
vzURLUkWS5wOUEno7QCY2BDqypKNV1+ZdDiHUv+sUfIoH1eBuMq25bWFJbLLVjN3
jTExpl/nJgDzeLBhpEM+ezgFJWZVB1m+rWuXRFbpbR3Q+X01wTw0adz3xcMHYQKh
RyZEJZUaNsvY+lSoB/3vjhMg5YaLTF61Xewtb/yO7S8bvgnYgKaVPaYE7QrKsr9J
/vR1iwmoglJtefP8bQq8L55m1J6AuvdnHZ/X5RCfUZXeMepMWxeOktfVnfXbcoXN
rgCXW7NR/4XKXCbwKvdCh1COuDXuTvdkhqxt9kPLFQNHE05KGj6gbQzD7xWyFHE5
AETCIktenigpZ22FOwN5BM3bSTWwzYY+aVzORl3/z7//Kr6791lr2BgacQviKHzk
ctx9NzB5MikxCZoXHd9QFL1eB2wpuFpj17VO9WyTPNyBk9X1yxqEx4yXw1wVcaHd
rg70bSpck7TgjNCih/7AYKz6Be6IvRFmGM8VPZnvFRdIe0djnIzs64NlzMwtO/ay
RjIswu4smnMGQZC1KDyedGZWFuDf7hnKoWYDrt20IiqRfFLVt0oNU5b9ez+Roc87
BLtnN7nlJh1urj3sy3AVhwZmys8I5rWuHnxYGj3ywKWrUtR5R402p0cnwPOEB4ex
TzwRKZ8mzlw/aR/HAibz7jsPCFE0aQxICnBqK+afmUR2p0g01yC2T5UTVo5+ui+U
nW3q1Y7hHtisTi/+D5SvhczRTtOCaSRRGwCjbMH6ubEpUzr5MrtM4JtftVgdAWPN
S5NeVRtK1+Dr7sdDlYyywuo4FORTRrgRdcNw6CX8Zi1M6UPY/g2p6HRrxexUK3b6
cwf566ZEwO+x0cIIk2KBd11ONuyFCfTCFmZC9TFCpOFwvkXOAz57zeW7Avn8IBkq
QmmjZDQJug227X7X0d9VZUL/7XLLLhU5tbwBqXkl3kv1r5R+hYVy8Mnfd5F4860K
mXJ4/4szRYzqpor94yuQ0Gb1r4VSQmxpIOv7Y7J5TRvUGt/KqF0OYKcjhSJR7rXG
vYFqsIwcqZZ7hY4IFcAs5kzyxwvh6NFQgFZ23bkK+CPcCMqAGL1d5a0GRQRRyBwJ
SumHlzqlTGJAobhlKAYoUPCpWTag2svzb5Mj07Vkmk5eV4V3oGEZz0xiZzc8r+YR
tXdvQ7cglZQwj6NIEq9z/rxOrdF1V22IHCOcpqSeOu8/dT6syepDG9v7QPN5gwVU
vehlpfQpWWNHOh3J3/zGN0IH7BfwmCR+eyDQie3yPd98GJI/VRdraUFRcaPKKtCH
qm1hbgaGXHun4b1Jqk/6gDek0cDcquMSFsRf+5wE0SBQSXjEMhd2rLETHKjOzH7v
8ktmeBtCKT0IPmTsq28BGVob8YzhgN7F+VL/wJ26r5AsXwe6S3x0+i2dIp7+GRyQ
/DBNsyaEl6khcXkxHI8JNwSkq8bfK1Bj0CPDmUjTdPUKAX3sK5qZsasd9BNh8Zmj
lO9MpEDiryr3KqS+Dm9cRJZlHfGFfq/tNLgJOKB5MpOfXLQx48tgAr5aak9JDbtP
VNUUZYSr/zhItBuT9AtTFHHBeiXVNCvxOfPCZfb3w1PNa2Qv6qAgpC9nNbeVaIkK
nNei1CumjPH9YXlrUukGKq82u1eoSDs3Knkjmdt/mPMzmKupvB+IdRfsxMxDX+gZ
ILki7UBQYl8uBzx1FbxsqwQJCagDVl33wJpVzyPBxc6ppbElL8+f514uM47tkWZz
w8c9hUIdLoyicVJ6/FJuCkLKO7attWdXiWpvKza5cQ7eUDuiWn37fkK7ToGbbIbc
VuGVz52k+OsxDBGQVVh/fWfs94gCHihwCMrbnnMDcCvPxhZ07K9a+tf0kCfO9Hvd
KAYOHpyNZgqQeEESNqTbrVzafJo0lQy5+sAwA5b/OzyQNvSYLQq+zVd3aLg5WKTq
mz4IeXauTqtJA/nP5pzBk9HskZfRX89lA3fo/boc+j8lCO4Q+1aGZ2yYiL0QLQeC
gICvTeoKoVDE653CrEI7Gwh6QuAhIi31BR0cyGfvj7ZJpWkHviU8aQIh3rrU1XUH
YRI+5j+XZqnDxYkSbyMKvmfXJLX7QDScPGfJm9xVie8X6xbUN4rzUATraZZE1b4G
I+fRUkVCp/pY1jvJIaMYvzGrz6FYSoKP/cAL/OMBMh6DBxAlrjVdUnVF91bSRHXz
MWlCT9qqUP3iwxbqGMj1pS9oRRKSzcqoHnO95gDM0vzesH7rzjUCdJQSH7KtWG/a
RWMKDriS8ARG3zMxnQdNdPzYSyj1C2cHTyz9rnrgxtjEllkANO0XFUHvdWtLnu/t
VlAj/aMQLtmia4J6VD2bGYC3KgjhRmLa74+JIY7DQe8v4flvymB9plRYo1Vmi26T
0NYI5MxHc4UO72pgXDqISnVe/96uoSllFBKFK52XudIRErGqdON6YRMPrN3NbPkw
XaeyUxvomjLV4QY9WOHm0n8RHxQyDsZBTe8HqVx0dFeFAnc8mCbqx96js1xnc6Fz
lgnPqOUFtkBL0sFMzcJ50NEz+Oi0xhrpGyifA2bj4Dy2IzCVuzqrSU3qSK/l2t5J
tIWg+sMFqJXMK60Emsu0PCWFcGZ2IoGPVyqTqU1FIY5DSFm/TCqN2zBoemsYa/45
5sPGxZNSIIBfbUITE0+69O1Nj+nTzxz9Xwr0AqMZ6Zr0gL6KGzXSen81vNd690qa
HbfIctQLPo0mgXX7GVBZpDclH726PpqKNt875UETA4ZGovR3rsOE1AzVlJjUgaqN
rSi5M7fc87IrMQ7yeGZ6swtP+DOWbuPOLLglrg4mV8EaXkFUYYMnUaBe2/wLd1ET
5kZoGTVGUae9uYx5pkSgjTBT3labY6aM2Sx/c3uJrV5IVJifjM1CiybK8z91B0kk
jaQUis0u5fZ9kPCgg1gP90/x+lyhfS4XO1ejHQvrMrAkWnHndJzE6aY9Vk/xrF9s
b2uV7bCKs0f/SdjQPs8MgxI+54wEhwnrr+w6hNJLExzh+oudtlDwcNMEsZgLxbTG
EWFCN6kwVUlBza9ZHaj4yOFwxJ25UIAsItoeXN8gNucHgrxAu4FKYnjR+u5vgyOo
Hh12lhMfLk1atMhtBmZgJudqpHL0A+D4DVjE50vLcGSBKr84sKwSVLPF7Z4KYbXH
JyE/cggQtXyzvkSBdsmymcVwasSC64GmsEVcwFTxqh49j47f2S0yunYxMkIcr+tF
XIsZw9g9V2zlaTBYbHCfwax1VtwNbrCeXHZrMIKcES91bvhBRJlkxed9CFRNpARU
7NN3+jGV7XCfoUHktFNuGdEx/KM77HsWTPB0jwOjWPNk0UgTtt3CBVnYZ3JOsIcB
Zj2hj8+89d8dlOdzfFruhpnKwGLqtF/sMXz+/Mfq7RtzFJeHifC12acAU2vUfPam
TN5Y9sh1ye97Y4fvFmhxyb/DsT4geLrvMigFK5H7aPj/gKRNV//bWnJ4CgWM++pj
8VhQSnRt0YyYyfT/KOGCkqi2TJQRG4Zz6NpB6XwpbyCjpXbEpDnJAviWIH+b1HFa
kQ0iBqduHGJYZqy4Vug6hXT13vh60F2bQeXtF9Zv7tNAzCHCKUVZJ/u55ZhDwGzF
U8BbKR5sCCJMvgbpGGd1pb+TSmUbJDySEgHOEtEoH5ffWongCL7uYpMdrGr/pSio
KZJDdvLCJuWca5/OHxzt7EmyjgHXfKj6ZT04/QpRdH6dxSABjyGVdzkEIYVx7u5+
7UjKVJEsvf0nXn9R0vgPKsN3VC1b85txEMqpENGWqZWldibmRoB1gu9BqSLhWIeK
vj61XqV9+IeKALsirE65qhsA1uSu3YCAEdrvEaywb/hC8lg0KtPZ2w9PwX2zcW0w
YEa4JxNc3ZWeDILB09lPtnC2ReHbQvsMttagS+sS03TB4Hk7Ls0/CnvKg30yHrxV
k+bCz83iMu1WU5cCwXuXuz/J3bdttoRie6gyUl6ZGxU1Ygd7f/4lCAeDYfwui/DF
dGI2/bO2aHl7g7j3zruMDuqBDeSN+DVaFhs3RjIHk1iwBLoE80gu2ZgzRu3AiIUe
fSPGpwXxp4e0DAmNPJTjIUsj4ZjCw6hdXhPiZVr8WKnnC9MtLQ5jONAnEKg0UJ3/
4JnXCmxXW19uehAxVfKNyoiufus/cFCYCv4tya3eduqmhnWbYsX80c9gxAxk2d3C
LrXLYd6K1ZcJcvz8HLr2RAHBRBZH7B8uG9HEjHEKsVX+AKuiwv0HKzZH3arHhXzj
WKXZ0AofHbgbT0T99wHmgurFKcXHMZknQKTnz8FKl9yb0lyPywcpEUzwVEv8tFMx
D+UNUP5epMertrsWBwRs3EkUYFj8DRxJta82c24HMeajZv09vONCPNliOq1sA0cf
l09aw1jjgvZkogzIR/JNhxK3+JDM4qnmwzFhi0AbdfKPCfExvjPH6OuZd+PQz8eX
8ySh1DI9vkR3NDT/QNRo0tCkmQMMRkfwG5hnj6cyh7+lG1peev7Nk6dmcme5nSc3
KQPQuSCuccRAqpTgm0s7b8R78a9VIJ7HrPAZUBDvb1vWzn88xMNYfbKNGMIqcyEo
BvcZy5ZPEdI/TiSnWYGXGA3wO0uV7cgGe8c2hPgxhHIOg3x5lwQRLr33fu4o9V4t
AJffnZKIsaiK2YrqUnXBthxSa/6aGxq6Ol0uKIcniN436cZskFjjLOz+NlJXsD4N
vSm3eRx157OzIrIcbumtK6J4k/0iQsipiBnKg1ii8H/+Cw+AT6WzXLzRuLZqy3p7
ConlCvdz/Dar39qa5NYaHmwoKj5Men8r18KxoU9XKDacLk3xzG62WXJSpyBmNZ8d
62F+fFZawR+P55zdFAjPLYccMkVvbW/zhJBmzb/pt6M9j4pZ9IJnLn0xiydxkEtD
N7ygf5iSFx5PCjaY/PLe9t24xTQRHdI7vVc3tyWDzLqG0ezZov1DJ7Z7fqlsEZMT
3dJBp/CNrMXmfaVqfXaKWR5NloGPtPiXlssa5gU6AEY55ABuJQ6hwFPWOCZ9JIUq
z2TIrPaUupAhGFZZql1pv3ok5clVk40lP6IqV+HP153JRYHIC7keVtEVrgXshR+Q
8FAepTtLPLs/DQcK12WP4gWo4rleKtdh7fHw9xtlPgyvnL/rwA85+OM823BHxeeF
tRdQSwgrIGPoCawjn6eTTPvO/d+9wUyNNeFXIQ+y+frN590DiUHdUR7MkX7iT2c5
0APssvpysJ9QaV/BzxLjeAzaDjqVLDxhYdp45TRaDnGHrpSE7yvuy37u6Cl4cUhA
hgrnh5ye2avJUJaVPpyKjYdZs/SP1x1tEaY3nfQJNdyNd7NA8Gvo09fv6GNRYcNF
xv7Popdf4CAbJagEqAgzbhJt8pGDwZDXUR+Y1n+NTn3fFBSj9oEQI724kXlVVDWg
kLaBM9R69D09PT2P7r7WVS3M8BqR+7Oxl1ovSCg8iIwTbOvq6zFUTHH7aXoWZGtP
RcYVJ0LUanvIhw9iz/fxU/MuCgIl96vrmoS/NsSDC/fZQAu0Z+9BCfi9ab6kJ637
BJWaBPZ2ty3OU5F7cPpsVH3EELw6TRyvfygzqdE6HfF6h+3ZtMKEtrlsG9sNj2Sj
ALOPuq1gkPIAfA4wsZxBh4eLStOdaWIegSfrGYyx+oEA1J9j+0GvopthBHZQ6tcJ
Z93XsjI5vU4/3Jy2tNK2huoLdUsdur/beoQJN+v0iQiGWZAQi/TFwwjxsWMiySVc
ZeKPZv56yp+rb0K3gec+0P85e1vKOjXtJcr4rRcxApHixZZvZvNw6C/NFo1JFXJy
3KEBOLuY13uDdiOfm2i+Vgu4nwY97lLERWb5YSOFZkfn6FD1kc7mr/nwNT+ohC8b
ubE8ZMv2fJVD1uXKttiIEtDLXCJK4dfclp/hQVYto+R4a+TNAsRQCp4DI/YE+u7x
XpH8bwETdESO/Frp0xjl9MpP71tvIgTomaOIAVSSah9rhoGe2yKvfDhYhsEdR1YI
nDOTTVVnsgdAy1BeAdIbgFdJiZZ9mJ+xHzulVMs7BH5kltL1JPcgAq8K5yy08DtI
nY9KYTtxGZohRXQv45Y4rLEGznkwOVsJYpHE1J64pavrtHafztnOviViG0xzrxi1
M0CkS/pycfaUCZ08BipOgVjowwrSedRlSc5v0ji0O7zxO68TWlbqru6tRxi7jlIa
7G8YH1/ZvI1dcRD4lhEaC0BdFu9/wKLrxJ0TJhvaow8QL38+erFov/D5XBzdNvOj
ywmwQp8kRTcSchlJQbiM+N6s09Sk6wpSis85aYt26HNERUAccCrJK+RBlI+KL8FQ
VnCD2Y/PHc8MUmg7eOAl8V2hjlPXaMfV0A07BdofbAVx187wStE+U8oee1ayCN+9
6jZvcR0SBBpcTRNm0uGSv1DDuAZuABlJpB8KjDr1ASBQWXCadPdvGbP4aten/vu3
f8qCave9BJmeA07Hk1hHPwvpIqCxzmnmO7F001scdDDiz2hjeLFvEiS+nfUnpIzt
OipAqlO/f0RtQyo9N6pIs/gZlikEzydAtao79HAhjrB4h7KMW3LtpHZKQcqDQ2PU
iZA2QdmuF5OBP/Q2ImaDGq7e0GgeyswXgnzgr+F8cjRZEDG0OmNDGuDULsv1lFWg
UzTMbB7mF2Q73iSe/eiJ0g3bZ4SyFK2LaWc8b2EbEsozhDyMBxyclQocbPwLQ3Gf
6l5iLmED4guMEXBliYd/KPb8F9j/REOrs16ozhFhkCfwKn+FluWzoNC3W5gyBhtd
bMjJVzk5hACn4pTaERrKrt7+scqwbqJkRg77d6JJRfYXHXQI/F0e0yeSRNN1F+Fo
RYh8ozQ3hu/B/GcmASIPSCgSm8DKYC7FeLkIZy2bxIB/EwYv1tAecCwCeECouwPc
m3hzVpqEQunZou34pd/40CaI6OVeY4of8BwSqxMnwVCtBE9UpAWaSR1Iu7MYtDjK
m7xuWTEf/4974FM+L6PDjAgtEH72e/U67o8gqjNpcu7bTPsK+fsoBTavk/l6HcQx
keH//iYizAQ9r5qVJXPZ90ptXspvFP1ky+nsyeKm81Yh5z3yPq/EWzuOsaKbrqJC
5gxG1T1Quv0W7Krkh1gaKDaiTpTswqvYgR4kNPC43oEcDyI13FwOFZPwEcghc9vk
r9rPoo42pznIDtxz1n29xVTJ+emv/DGEmnJ1tnMl/ci4y5YVKL05Mlz0gsFL1Ove
LZlk2moccY2xPcdGrgdWlQ2le+YRTXGJU+q8kJu6VAhKKxXZGUjav8UJgcc75gOq
5u96WU0nb+b9QWf5Fr4cEbEH1j3F1y/AxbXeKtQUmG0Ub3KtuUZl8Nrtb/zADfeR
s++O0nf/9PYSC4iKFCNziI3KL5E1TguES4VQlfsp91s81lMPWudbYgIqF8iENp3C
h+dxwjzzRSG6upudNbBz1DH/rvQGmQEU8FAY3g3F7oIteEGQgvFT6DN8L0oRm7CT
kSvKF4bFGx/gxbcSliFRvqbDZmM+hQxGfIkKoZ6W8AzEs0bZhWe5CS3gHOrkYf3f
jB60kc6wPVB9FtA9nonItTjSbuVPZ2JRDITO9gnteCOO++vOP1JnskUgfR9yMRrJ
tOxgwtEHIwM4F/izB9+3J4xFRTdhajeHyVNAyGjeNOMTHSOKVINnYX67bGl5Ck5u
qt2H51jzgnb3ZxAyhd1dD84WpAB3IbNulEUn4f2K7WCvvRni2OJYSY/XEaiiP21s
uCIlLKvI6zjVce2BhEKN6UJxhUOKEgtUQYpXsGTWAu6CGitgfhyk/Ex8zugRX/XN
gPclm4IkjSU/BnEXwrDRRcRb+Z3xNnWVM8JzEXp3eMOi4ZZDwpQsB5uJ3wJf4QtN
mGRaf+pBrLrjOp43QUOgklOxNEW/2nTVk595yt3G2N/sJB0Ya03Xd47ZX6InhaZQ
BD7EOhI9Z5LdjojbfDrfYub4L/YC7ZyoYZTuujW45J0+9mA8c3+FMR1JAhClvhra
S/n0n5Vq1rTyyj/7GA9yVZ8bs8ZbASnY4Glnm+yJN1Vai3bM0qo/hJApycAGKX1s
LM/6cxBCgatTs3Grsl0NrlPzjF3rFvhkTKixUrZs1GQuwDBSMPcy8MIowVHMppQj
zPwxc0hrk5o+fOp+XIu8+906RACHMYkDCuMVnnctEp7cqxXCcx1K3qwBvmWYVrNW
mpjDNwnRWcdihW0nnqoWNi1/+G0NxaumzCEr+j87nbTyVMWPU5LUjq0FuPk8xvLe
zcbor5C9p9/nJinKAfTY6W+J89nDEaqgpK+MjUEa/CQR373B/gIipYSskfUKIlno
fmAMorOSQrwTFJ/mXfTzEwxYaJ3K0veb9iBye0ts94J4CLVzBUb7R+Vt2vPBvFPh
anKssHJ4aXgYkpJioR1z6EFc7oBia5BvJLPCrkXKPTlcSt9SoEk+MJZ/oANBajyJ
G5IeBynFGTHCe1U+QN3gwNSPJ/9su2E3SlfTyuAqY6Rds79zwp+9QfJiOTC23WXw
XE7vnxpIlarMYllc8QDbH/eJ2vp5fD/Q92G2ubg/J1tjimpmi8TcAadTk8DAu6QM
C1Ouob5w3bbWnAqwZ4aRoEmnQo2cLnn7EgpT4Uk2IHvwaTfne2EUpSKOSJ5Eqfxt
Otki2+ZvZfbGXUlwc0C5LiPRk1ZY4tPf7Gwq293s0Z/cYb0sBJ0v3YB/RlXG736w
9ALQPWkJN5Efg05sofZLVY2440Vbpt6Ollpxr2wVE38Gs97C9+K53Oh/G1Vad2PQ
MX2T5os89MB4VVYr+lPfIbmOHAmZrOlU/mluwrUFBDiFGBWfDCXnJ7/02K0p5JbF
njK/aItMZ5zCa4vJ2SQd5oZyP4Z8w/7P279M4V5yX8kfUfYtEucdI99zgjcKp/b8
Bp4MohIT96q4nrHKCcPND6EqCDeBbPrTUnIT5EBRexk3J5FaNDRBrFdB2/319csr
R8kq/HYTGnEvegSslnRVHOulrTaURscsrg6NyZ4jtTMDpygZ+yZjbhL3Oidpfh89
Zxd/9xrrjKpzUvXegc0Q6DG57iYaaVCrD79+bi/ttlo/oGUKI+lqXsATBv2LDdFC
VB3vEF2/Swf3nK7ZUMqxv5P40xmpQkY+tv8uywGj4jtBK1xW0eUBR9IQ1ThHv/dh
rbrUxXFR64S747LurBOF+FziNjaht8LIdBUTpYpf2qXTNGvXcUmOvd29mJeaoYTh
14d+Y8TvQj3qk12R69eVe7L/VnVlWjEP49LMtnFNQN7tQi7wciBU9M/AaGq+OPnj
8D0bBJo47HxQAcWsd0U11zFoPbyvtX68V0XurB3tJFCmhgVgAdse0+YePqqRaZyP
9aR2le3FZwjwb1fsdOqsjzSwG9M8eQkM6L+pz6ohszqXWC4vYhg+/f9BkhCoLImm
0V0++k73YBzcNnDilOcuYH89LO1A7O5Bvc7NKgMvwUAjbCSRles1Ls5aAvNcFKGt
L3RuK0/uaxeBjL/k4M2CgpnYqUkkA9ZiWJXdKkZKRu2HBAoGIuBS65Y0p3m5w8NS
XyJ9tQNEVGJJ9gMbMA2DQ66kt/djEQPtyLw6Xe7CdGmWBwNEsQyRMtnVhSgvopcO
ih47+n5o8wHFI+/VgioeN/ypaq9yY3IpNOMSxDigFoF2nizusDFyAgNUdKWBBT/u
2Kl5NwQVjjAmCaFvM/Z0c5B33Q8xEPm9CeTuB4/e1+v1Rfmd/smGcZiAAexlTWA1
39gRWC05rsVTXsn3hdOnlbcYY4+WdE827wnbFOyNQ4pnfCRFmQjwJNbubmpW54nC
ybt7gbidVSh6P/IET6keMQNXo6s3JWm3Zlq5iRVncf/bqGtm/E1BTfxvvpJBmC2w
R5f7VYTD+DJz1ZFNw1elPlNwoEonUpMgHo8v7pVBRSyzQg3Z5q5h19Z4PeNtL70M
dwsU2mZbzhLRfsC2fxEyNp7GGP0qIRUDvhQHOuvLUJ7b8lv8k3y8IkRQOvN3ztlo
KJsPnrboXTOXUexRPnXIPs7EvfzTIHyUzDo5Yxd7tTIPoii2vIsoM0yIfzJFG0Jg
NDC2EcHfDrSfuEs33GDodSB0SzphzBIQzhRQ84L7kZ/FHTC//8BvCfcl5OgaJ5oW
+Xf2idwRXanlIDlxMXdd5OWTUayWAB78XZpALSjA2eo05pYM1wY4CNihxFKa4kSk
r6mEYhzC2WNfON0fkePngL1Wn8HsXTfbBUjaLHUYmokAr0IP41jImd6L7EZLsLig
/QvtJUI4xC44XFjdLSRtBMWMl3xXNGUsvy1XaQSc2UMnqhQTFbSmZUNpSF35YKgM
h5XebctlOB25vz9vXVlffCAMJPnnM0g5dQUUY3BKOS6xL/+kYyF80zu3lNMYW184
mW6LS8jbAl9+Jhh4O7oLxK9RvRS1YFX5+kAiYi/yIAcCFkpsifllSPGhAhKHW5gP
pBFe411ho4cF1XPoD3Iw7YZweLHWvk3agESMHh3Hl45UmznNjWaT/vCnZfXzICNp
PApSIVVSUb87NXCnTdIrUK5KyNPbMhZ4E1ORqhmqJDE2yW2bE7ZSQdMWrdMYHqod
I9NDfi+vEJ40bBGfUxQRsb3wTkmOAeG9oyQdWRP6ATuvMXUz18B/zcJuPCESr6kg
9Lve12jXLdHbN6WvyjDVgYmixXaNe6j6ZnsO/BtZVyLUFaJypbVoLECYl+G8hmfS
bBLGH3JjL5aPw1Wf7NeTVKQQEFcLlGo+NoG/qZc4WHzkn5Wyhr7bCdgpbWkkoTLg
Bxr43QkOYcdqhh2j8Iug/oWLtEsWRzcCN39kVD1qcJs+9QcvHgb9ZHygoisXEBIo
DTttzgXBxKvX4OTYGdXLp+IzEPHZ0ruseCqSO7ZauvUeZbJm7H9yCgKc6q9Di2XV
mIjDRsWXe3PX1wVk+X/bd81W9byInIZdCbYZzdiM6XVUbyDIbMDHP1MTDsayyu0H
4ofEq0+BCnpPnj7frsCiCR1ySqr3lruM/Zlk9urpNBeKlLnO9xOsasfMA/IRolfO
lAncxEd415MkpJn/gcML7j6pX053bwnIn934ILq6kc/IlAzqeJ/Cboi6CkZBUkl2
uYP2JlcuTcg0foe+JFPegLamCHm3Bkd1S7E5qFkw+KbWt3IVhj+RrncAI7IBEswc
2tDs14UkloioNAyEY/EJ+d1YvQZEOM4YYUU6vaQtuCVZ8mLO0Tt2cRfNMBWy2jwK
65vmiDUqEkTp7wFj58XQWsx3ilPFvVzNJe65e5iU+4OyQZYeFKiVrqZs1f+CIAXL
RXtenm1HBFHpJBRwTdUpOm3bj3wJwf92PtpNtGw8PqWkmXl4jQrNCRH1N/FzgpKc
tvKIrVeO7fNhdbgVLwzclUzNctnQ9za7gTP0aeekCUze4Wc0D4tTTCPA1zvgjE3+
mUVf2ff/yjr9a3h++tOmNzsoW/Idd0Vj0P0/enUmbc0MlkOMP4l/vj5P6H1PplVP
W9uTPGeviTbKgxnog7Dv8BtbRfpzfEq//f+2hkYerVA8k5r22LGl7XBQK2lIMlo/
PAn1RSLDdPScWB6yK0UVsyhJv9Io/oxUI5zKrX+sxeuRQBW0TcTqAIz2TaihZivg
KBQ/MVD19rJX2jhyuDPTo0tL88sA1K59kQf4V8/3NeWD+WI0Tp/LHhQcA+PpJGLV
J4jF+7tWEa6p+NFrFwhHpdieSVav6nXDWIg/i4YZRO8+UkUX5DehrpY5f/QmjG6I
rRJ/9JzX8eiZYIVzY8TKENOS2X9aAz/7vKvQTn/ENIoxXE6xXL/sg5GNbsufY7yg
ygSEZ0EVuX6dCGc68s4K407fVAjZnLKJ19i8CtKyQ+ECHwSGrL94EpZLMPd/UnQQ
2r/wT0Msr1Bufc1oYcrQIW8pLvhj24edC59u5eYjeA11irWDiE2T2T7waIuBzaqE
caa8ScXQlZeYswqNLCxOh6sqQUtTN5Xdlm31sG4PjPlnHbAeGQAzVuYAyynn4pJe
k81c8CpOlHoVw70gITwlK6X1id8zU1aMqxaReR7Zbm5tdUf8qBySDzKhfKNMejMS
8db0cWWabtERCqw2H5WYwKE2kSF4XqZwt0t2SfHGlJLUFX68rXRhR3pFpmoltqcF
WXqaJSRSnJMqHqTLV6G6hXSop7PJ9q3DgZcIp9GEzvbmiJwkQ4h4m/qKYbJ03cpI
uTUkgianUchEiDVPbHyPAxoFvXgvkpRt9ZtaYCJvBzfluw0ZKKoJlM7vPzCGmu/7
fG2HXWq97Biuzyf8IbSKMo5b1beIL025Tml9KrvYBNwlq9uQ1vZckG/zz0Pdk212
r0p2stzx3Bq6S7R6KIGjDUlMzqVRrCDHAKrbCu2Z5eRN24MElP22lA9TxVpnV+lg
qGS6pLOetCFLHGGwrTZb6TlQBHR98Gqr8R6yO6sCMjxW7CExl0zmCzWtHg2+3uwg
Vn8UKgg6oUQJ3Y7tj4k7wkAcnx6lzQ0Cm0T+AFhQHRND0CIVlSQ0KfWrK+cTSYdD
9zmLg8IbVFd7gZeVltWz/veAFKvhW6eNqGNBhMMClEE9yCuNf3WfMgckzFv+Puqd
wJqFfiFUqGzarV6JeCi5YwTrctcgMEbxHht/kdkaqISxbGH8nm9CK/Oj8CzxKZTi
xi2FG5RKbnZPy+yChGa4eY3BjVo5YJtBgu/H6fYRcqIowzqCR/X1lFdh/j8U61Mp
8QJEwxdxsE2JPCHZsQCALDQG/YMwX5dn5fieIyZojgSytDSCkrwaWYpi8wNtYomj
ZfHUEBMpq8c/FGlYojLfzKEng43c7PwZz+szoe/2XgpvN5oPiTBh+dGj7v93KJp5
/yIF9TqAsFoTWBucYtqdGOKKUBHBQovmBIPAfo961ofNlw8bZ5ipW+ofopIimNST
gzljug8yndvCFZnzKiZYuEDcBkVJoTZAglGCikklGW+XKTtMxlNp1ganuG/vuiaI
I7zmOhYXgnCNU0m37fQHFOkSTYqp/TEmAy8JYEUvitOtvl6PzD/XTlNta3HKCmHI
jZ48F0Pw1U13HQBticd1Z/AurCM7JDQjgw9lMrnT2G3lOlbIHP36DFlYuN6Oo0i3
Vo2ha46U4FkXnriB4JJzCAYif9d8qcfgWllxR6BTsCgT6ANS+Is701RRwFzrt/1/
2eeOlvuVAfFMBNLE4lEDU33tPBkbZ6CXvrdPk5OO2k7Gj8YPGvZhtX3B9z38H3Sq
Aq81QE0JtRtHGx7cm5/RV4fPSYwDslKj1WOqLKXWEwiK6iWWQTRwA38ajsY6747d
5msXBCY0kNpy9y4O7QRTkGF7p+6hucWCjhZpq/GAGThXtax9tzwvIFg2/3FLcoW5
6isd/xa6b88zjclCQvJRj6CYc6FTIe0e+dBjeL3XrXgQIi3gF11WG/VEYIVM7M4H
S3/BePC4/YKS7/bpkjhdYxZwqdKNO/0XAVkRDxWkHFKBD26f6od0YS2Wo7WL8iQE
Dmx/OKYB354uPfIBxxLcrglPOQJpwyiUHm4pWcX6LSETqOKTqVmzyunsKMyuqq/d
4TyrQ5ADix0t5bCF7oCg6g37Ng8fwOBW8EYRjJALlpY7nqIHJZqdJL/Eyn0T2FGb
DPsZklgn9I/9Q9BDkWdo9S0x8LTe9O1xmpA47avjJWmuoDe/AGoFgCWovbOP1wmT
rMnGPzpIH19x6ACnKKmBG8hT/TGxjDxbRMHTzIaNQHGNL5A1WLpf3DXjAEyxZoLK
rg7C+bsRmpkTDl0uqyLxbTJpmnKm7v+/9K6KlizBeh0lKdzQKlSPQfdO5I/WdYrw
4ibcDVhokQoahWrHFgv+dr71AhYk5zr5+aWn2BaaXjAhJitAL54gGiSoP1LP1LYv
RB1/PEAOUlH2De+XnpVOLpoin/VdQG7Xab+pOiaLfmsrVNDUQn7km2NFl5P3iCU0
EtrtsrY6/5W5rsSZokD147ZWJpJ/aGRlJSJPFbtmL7bSIyVIsoW2nHydYAV4EZxL
A0GINvYFaXXpmdGscYp5JFCUzbBkql24bSPa94ffIGp4J8t5llZobtEqNVj7RSGJ
uE6GRffx6LSPng+892ph0xyeLjNeR1OyDp9YguzbTyxdieNOEhwvdu9gMBRMEedP
KA7tYIAwr2MrM7ifjYDVdZVngvAdfJJWnzLUufNm9Mbv1Dup/A9bzxq4aXJwEpKM
KKdlre5/FelGr6kvV6ruHHIxEWzVWRe+2RxzJT8XSGmsVvleEVfTHCKikXbxMgqR
GBkLSOVMFNmMjh4nxHXoWQvKlxv6sD/XXtgFcPjjeI9V0K/jMTI5eqI8RwOiplvf
JTpM32Gf9NUGD9VwP/aMtL29tXc96daquXLIYKrqim3ZrIYtFZRw2kak7lYiZ6sv
4g0nm8QoyuUfu9JEiKhOQ/8J4jJpzik++0aRoQJntsfQ+G9LN8h4oarDAoXrQX6t
CLGiZYmmdTF1zJ1KSs8j7jlN7mmiKKEBUh5PQdCB3YPdebpTmPDracki5+toBEav
uPvfMdf72IuYJPFJysimvuEwOib2BEx78SOOGexp2zUAqJJYt6T5b8GBpO4EY91Q
FnT1oIH8ukYU9yZh7dZNjvFDuSuoqUOKgXl5bJs9WKdcW/2Iut/nqNnFoD5yzXYR
G1H/UCYWgMM4KjGxp3k+3NRizvOCcaNYDYR80orwmVZJ5Y9JcX0jXmZ2wtq4444g
GwIjl15Ot2eIX1FLQZMnxZFO0FmNyZ2VT2XUZIOlPJToePhbSdCMAgI+f7Dm2c8X
/oba9HjxnehQzA6PoDUup4aSfnWAyxHvN1k81P0B4E9ZqwiKHyGZADt9mLdXpf6R
Yw3bU794GReft9PoN46TavUrQZ9LqZ2st+UI3vbW+2F2fDyroBcKalzpQ1S+9QUZ
k9XmxZL2HFi64SAPILOt49+G5UhqxUDpc8jfzz7XQs+hbP74ZEqO6Bg8aiSFj6cz
PpmAcqBM4Ky/2Hbxg80fdDDpuN7wCk22deGw78R30YqOxeM5v6xll4adOcJ1Jm2u
QbYcUP7uUzKS+NimjzsvP+BmAujqqOv2pvt+PzMF+dvZSWMfNW/Lf4Tn24s9OjWd
UVea7AXBQeO9BxyhMDPZXISgttismXcP1q75bqdNl6cRvX8a/ZHyVuDhuyz1Mq+z
tsOWePd4fXtszQCNQ4im+cRutAM7aL6xDJRcFKN6HMexrHRi/8QJ2DO3alBxEKe8
3gcmgs5klKgnJ+4Rtuvj+aalqVkYlLyPCGgxV3dAqbvV28uLJKxewpN2fkE6divz
2bRXthNxl73WVuGYfgRzYGQqxYgAwOUwLXntmQou7zYX/QdBVMHl383R7KKh0vgl
ddQEodOZHAz+acKd5tGYDcyoBGDTroB735VDFhHWneJhx0b0lISrp2XSCLdIYCiS
1JNOHsm0U+gncR13SzjjoFx36AujztoY61mCf2w5TvfYiiKEDG4ksacwdDsMTNbs
iB0V4ONvX3OhOl+2EyJn2rbbj9rbEitcaBEyUphZZvosTx3Uzcn2CUmN5r2J9moE
lPGOrs6dAOgAmxbOQAWpywXT7EYGzJ2ReBvohHDBolt8GffoTUKT8RY7nPxjJLis
F84LHd9UePYi/Qxa22uCCOaUksiw7QSHfLBhqr9bDYrkC7UDU+J436gOP7nbc4/0
xPPhtstU9kk3Vm/+iPf2bZtLQ5tHUQMwH4J5cYiWtnKhKI9QLCOjiviv2yg5Hmia
epne4ph4fydBieINwoYjwaCXiRFztlqND7UC5kQX4G1tcghx+l6isW3zRkdprczw
zPOCfRHcJ2vdEN5haYTSlMW3UMH26FZe8tyGiIQuzoLQXO+D8oLNLBqAW1OdZRqX
vFii1ZXRLad1HhOHQFzZViLESOkxp1OhwSLm5zH9CmF+zRjz2ohhQ1DDTGp4ZTfN
r7FcdB8J5e4ohdvgyb0jXCwL1PYRz6luQo/tsfJ6fga2ByKJyCeWEsqDlWF5Mp90
XO+FHBqK16MqLdxg2GCe2AdcklZkwF5dAZ4o74eZlPWD2CFSNOvqB1NqgBZfvEZo
97vm5Czxgeivt/3Oymlw20Y5P2erBDKnhukgSMTN4TwLc9KEY38jXGbI/amEzDsd
RbjI8N7MRoKIr/gVkq0HEA2H51EhQWaWxoP8tr4JP2JYNUZGkrk4G3gLkRW0aEqx
P9t7E5sMU6vS4TeGOrvHXNxqbc+6fmklqyKrsL0LODnyPOzd04ha5mVF6SwTj+WH
PJncGRCIcC9IZkOMUkzyxJ7/+RC/7Wp0iJjP7z5c5oKvNE7CZYDhqKO68JO4MVmV
F36MM7QEPcIc9uVPsCdGrM+PetoEhCYjA4GpVNvjr3i0ny1zsJbM1yIQntAYPh1E
nFx/NveTH4xTPeSqEQbjL0C1rSxYWZE61WEeNmHqVKO8Zz13nnBtv0i7YFVzE22d
y6BeoJhFkI5t/+c7q+0JnuIkPD0ZrXkmu79k3R+xJCc0iA2jwfhGQKFbK29HeIto
YrwpGTwpeC9wdEqZcByGPV4eTxAhDUoGp3gp7VLdOBzImTwepNKn5k1Kj+7pdjPq
qZYfNSWOX+722YSidPeUgQGWhqziFLczPjWdTkFAH/Tj6FRpZmjPrbvGF5zO0Jix
pk6VU6xVQNkjbfGaT/E0eTNtJN+dCD1iih0kHfLGKrMV3xPM7j+zeUA32Ohc+qhM
ElLidAzh4zsSmpitF2KQk5T1ugSj3nLbXFTWoiqX9p8B7MPbN6yiImqnW7nu90Ho
gs2z50reoQJEpzqBYQZAtrsfSXp4OHuT3bu+ckm+Of0aNTdgQP4EFzXHtltypXrV
mQl1rK1VcPDceiWAJztLjefThYPP/6Jf3SgfZ/FN2PINeFGIyEBEj6NUoFkk4Dyf
6Q8dLOcVB2szA+FIBEVK5t8zQD/S51RfC95O2+5nF1Vqvfe0Ti/n2ad2GyKRtrhY
d6wkHwmvg2BxXLHe9hFSgF562ZfFA5B0aasaQgiPcgWXN023sdl65lJU+s2XBEww
U4oBxHpCaAc5r4l3IiHki8VUzaRfi30xJJBMCGxWTzrNq/m3fJqbpHyd7HX0MtHT
v3IEYG+SaNY+I9hCNz+gaiPZbcPs+mSDLWgz0PAZwSdAKlIYf2jstBE1997ud4k2
DGGdDosDGC+LhkGy/3fjjLoNs3pqve87jN5+kHoiPQrwBfW2y9OhTLg4gQak+l6Q
2ufaQVFlqy5jg3nC5j+/PJlnS3rYU5ild1uwk98SchMAuNJxpBDLbgOly3Wuozja
zVpuoPe0hemV/DPrUHn7ULAEu/dQ8eVe1oIXWg/kCuei+mObTSvdyoZpiXCfgcOg
k2ok5fZEN/qJ0OllBGBXPZFu4s8Frht2R0JY57TV1PGooK6P0UlJZUNDgCLW/ZPu
MINjXtj0mjAeNgyunOGl2nQaSUxameM4rCE1QToA8MV6lh+lGPzhFaRY+Ik30aSe
oSEMwCeafamPS2aSZTnVZOKKG5jYcmYVlrwBBbhGA2IooC1p5Al+BLWiujQdsP+V
gGCX1CdkqR+H0/WVoQCSsykOacHbI8Kqu3azwXGtWwxxew/ieCNbJMdakHv1QqbZ
3UUOp+4s+MAOsptKONf/HI70gFNvo08HkM0CrGRRRSbyHASH5ulLLUSuH26/RW/B
PY4MH4mJ5SpwtTg7WJK3lByXvRzd0tr+bwIl8wwQ6YyxYEF874iafZlhH++wcK8j
qvAuInkJ4YRfuINID1wUSAv4kfJCr4IbmRuED8ICgPwHy6pUmRijCukeDAFeEqlz
IUm1rHV/hwzSNUAl9tOIQ6FyE+QyCKqQPzSOYdN8XnuElo2Oh1Gfbj8fAUTK33mm
gzgl2J/t+dJeRWIz4/Gt4aQ1Ru8ALxR7ByGSbs1uqokc2L9UaRzLZdIs17+4pP+X
yI5KFVAHacQcBwJIWbq22SJzkdMMBBR38dIE3HeLzRtx6G0ChK/h0+TEYHhPEpuH
ooqdARS3ykVsKyf+xWOKJscIhoR3m126cq6QZsfxcyCI8bRl7Mqvrw56Hxme7x/F
hII1u4qwss0CLqPVEtxKIK/59tM1QGNKiEhrkTPnMRaBNYRtwdGD7K655mXiC8Nn
k4Z0iWMdU7E2RV3BM+GOWwLShsni+TA0ELTq6pu1hahAcGzeo+5Ii9BYLAnOikzf
lKtATBV6wQrHdwlsCDAbFu0wsJxpKR2lbqnyXgsg1agSHMkNKcOdtdnvCuFH+XVk
YtlzNH7yxw1Pc63rzioKo6p6LrdlJOotrccllbkpkIv6YdWc47AZuSKic+Ue+TH9
cn5zbPd8mnyFL27nhCoDD9fHywVQpLUGPWTb/KZ4zXi7EjXAWqsjl88whR0QXQar
HNi3e1z2YGnHFTtuG26AoPRc1zrdh3TmrQTHbK/LczXbj2Tr/iw3piq0+QMZ2b/O
eDnFZvpDNSjS7kJRTELtp3Tm1cUZnw0zoiWVUq94UO7Lb1zA1LxHzks0cZ/iAHgE
+1UOjCLFl/LUxlftBcwtQzvi0zf7vCQ1DnwpLfvkfEYHIIRxf2Gi+fKQjawWZ897
rFv1g5SBit9S1aTVJtKxtuLCmc07+/4ty+2dpjs9kUNBooOaj0BY1WLfE9KVLB7V
IHZRkrHxKQZvx7CwoklwMUeZu80I0jYGzrTtSACwuveCd9nhEO4Dh4wOXTNkQp7P
ovDxYPW5FjMdrzVJzcMlHZzRgHgL8hsKtfR0PMvm1XLanKkXEExbWkzhPOd4DRna
Qscu2KA818lBsszxoNM3EbpT9PMGAFcGQw4sm7ryzG1dPeDFAhddhCmPdhyGLJTt
UQPpWjAzoGEbaN9AGZhZaKFzR9cOSFTEtFDmJ9aIXQ7VbxNIKm0okitltEnIPfCz
3Lbtr+CNYc3fw7eeg3l0BHiJ1IZRuK+mFSEwvNerRQgGlPH7NpFrsxB0bWL9VDGO
1QnzRBHGWX6BKmo7KR1u2HaZJklq0FmrBU2DtPc1TdRud/dkQDL4sna8E38IH0rd
DazOCVUZq3YR5ilzDg1Ox+j0cbMBig/XUx8a+xo0nkTQIEczfawI4MMkmUDC/or5
MebqnM2l7C4VHrIiXDLnLkxPqDVSqH9cbcYxkMBZfm5Ku10oBEAWPZLJcTP4wIvW
UHZhSb7CKwHrZ5e3Ml+SQif0i2jbXv7wLh9B7IShE8pIOC/noIpkhvjOD+sdFPUU
7nosPofmqVY/n21fcBeFsZphYJ8Qo7WBBvBH+/fM7Q33hI+yqnoh5jlVCIMlvz5g
egfxG6ponvoQaTk3adqkl9z0sCuAA5kuxQbhP5CV8mDT6kTtsQtkbngoZ9gJqF/j
T1lN0PKUZw5nkbcDTGRVazmnKle4kBSmwAwXYDEzrxQwnlgXYKYq4HxL7rU6KqCz
oN5s0gvK3QS/tZV1rVimS8LtdPDQfQBE98TQWk5sHgZtmD2Qp+YvXt5xTCFxVgJz
nO0aWvIecRvpXJijwMEteLTknvUG0Sbwy82bsv9+514EZg2orl+JELRcbw8LRImm
Am0rYQQmWj5ZLqiVlvBgwuR4eOUjEHCya5kfqJsojU58uLcSvnFe6WE7+AfBc47S
yRZhXByH5np5PTmA1U4YA73REjQKt8b6rML5UmE3+5coVs2udilwAnEoXPHo5l4G
eVmdAaNoSZVfy1o83pVT/9ZCWcOnF0yezVFhWjOKltECVFP5JQiUuLdayzJ0d1sF
NF+Q2ETYyYe9LLf14PDyeuX6W0zjhnN2To9/OByznWSZQCYOsQuGOCLC1AP7NGtI
tOqoQ/2vv8y1n38LoqGnkZTBpSQzYm3F8GBxAmX12BnB9UqdoL7QhFdF2cgiY9s4
l6zxMTdAWp1kN1ZdkpJTQiX7iptyuWY/sPhrFwDvr46d6hIBPUBG7gCGXNL4WU84
n8bZWRD+GceDQlzTGzFZCgniJEZGXrgV0zXlPR6ULWlR+SVH+e5gayH0y5Gjho/k
IhxDM5SRswLR9bnu5/rzRMOtQY1G4Rlq/as0DBFmOGyDrhP9akwYqVQQpJTfDj+j
7oMlV5y506JPLhwkcoXE9a9MKLes4pAoqKp+iSfyALmjtY6pCI3VwfLbn92MI/c7
XSBp6e/zzSgi1qcNF9WorDrjIChAUVrq62iP1iX5bHXKitM7VkZ4Th0iIm7mO4y/
tNGBmFqSn2qmTGMq7K97Hh5yy6BPjRL5eRB2fF48g5kd1d+PE9M684jYfswY8yYQ
H0tert4ugWORMxem+8B8gHK+9s3xXdBhSnue4vH53zdqsL2ddLfdSlOgjZ1kFHsg
ytkxy78Q7+J+lnaJAjUT+EeJpKweMIuPtzA5JbF56gnLvNhnXVfMgHYubxvgFpJQ
FnMQgCFwHbYv4pzw6yW61HRktp9IqRVEsTYqNFoVrZ50HcEKVpPqnQ3roRubYHjx
fJTcB0TO2M0L0eiMyqDjToJ+FhPVavzM1wZMCp54lJXDzO/vxndMyY9/csExUsAo
wP4ImpYuAeUDbmh+t5oGa3a7a3N7sngcvAIsq+8JFgZ7pN/wedJd70fbsD+Dq+oa
jk6XvOTkWOVt4/IUm57ISQLVA/09Vivt6jzZ5DZcBVOYZrmNXv3qB4M9+etaxSO8
1tLkJXUJeWIEohL5/ehGG/NoBIM7Q53yb7MaNlIok3MBJ46ru1Cz5VveQJ5adwrM
vUKL4VxzqWHk3hAB3P8RPH7Ihz4SqKbj6niz4AhZ25tFPqJoDs/UQg4f0ierkxs4
a10EopJQ6u1vHSuxxG4w8bYw0J8Ima4a8Ip/ZB10AhzisvItnPFAbYB0HdPf0h8q
JazXiLET5rSjCL2THom8BZcvjy8XcQHuGEHqUTHbnONb5aVHKrqF+5oXSt2u7ALW
6GNSOj58c2QdPyOnoood7Y79KKlLvA78Pm7IuzZNvbSbjIF9WZsxv520ctrYkFOX
nAu3eagbYc7/LZWhpdWG4WNII6vM0/os7U/hzs2xo+XexufdygX5BZRc7SiqekZy
zlE42OFp0ytWiJMLepEvw7d78SyIE/oIO6t09G/ETfqKhi8cphJ8/v8A3l3KMYtg
qRwBKaOBruzCoN4ZFRABN4sqNPwO9Nn23ILOrTBSh88b1zKwDgWY2U42mGyVbGY7
AiPUTQmumjRdJT00voUnAH0fBXk9iyhwAogDuuHbMEgIoY8Atar6Joqc8C0YmXbS
SnpAa2lcY33Z1r6xQarlz8Ih8C6I7ceaXjJf7F+uNHOf9WVeoR0sVgvfn4d9Dc6+
S4sKYYyCKQaC8a74wnq6lHod9QnZ7IJFuFuvJbwGGsvba5bhj13VBX4h9XUGF36l
ndXeX9nBn3k39u5/E6nHXrUx5tKiE20s3AE+e8mhU1Sg76+HZMxIbhoBuyWY8333
ALFhfbHbIb/btQNUonKm22SEuL0SG+1k34kvlvGGKMOOdPpLMkHL8ZcXynOBPo/K
TzuO7CBeMaxfmgT6WYzb5wOkSnKcVF8jKKhv0PuOZKLXoLksGBqWRxdW7w0XNHmB
TDVONW8O3zqYzZpkgieKuO5xu7IBfzbvAe3HWN8RvjY3Y0sEtjaCjsvK5mu9QZ/a
hNM3kCWVp9QvOu1WtQluMnGL5EQj5kE8NG2drqn6D2D/3YGYCkvNVWLhQ6/iyih3
egPZsnw9hxt/X1DiF5BF0tSwaEDhNwByeFjaVtt7nqQzRTnORJHnN/mSOJzeY/NS
A5Qwz7UpHkHed6R7U9D6IcfWSyYBL7yF+3wxFndjGf1A7m00wOGhFfX/5GzxCaPY
jNuPRva7OjZV655fDsGtvwhfQLpmxrgvC7nA4+Mj4ahAeuBNNRnndTPf/+SR8S+c
DB/LpiGyqbWAa4JCvx1UBtb1hww8X1eecXs0V8luGAM//oLsBLTt0yhJTcbpJWwn
RQPjBvLQOPnBjspAsksjrvZfIGy20Sl4xH23mwcvRkRw1wLgRwpEaEQ3yfZqoLXN
NPKBzXiiZS98wjmuggwfyYxeDMMsRAWaJBYmQo23E4iPmmlN92xv6SL1cDaaqQYM
II82HRMxKXZD7JSMEnl3EYfUo5SQHO3BqvvLmbuFm/77xj2fH/gWQRKqH8wdt6TS
v/7zQ2+HONLAn1w3a2HjjO1iP8GKKSu6Kehs8ZW2k1eu9KQwq7HxLtLffdsti5Mo
1Zh+v9HD9t+xeYKV6pbED4roTXJqTsj/O+uRdltaUr4cljeEZDfTaTOJD9qaIfEk
PoFBciEuvEDKIBzyd2x8pcdzxIl+qrAcbRyXo4syWyYjog25YiRZ28Puwi8vVT2z
YEamFkoCizHdGStLeaNsGCvTejs5tRyGnQGholIOA4pvLIVI9pKa6w+4euMu4MGR
hO/heVQpFQgyfvdZfA7fo6e24eDD1LCq3+pwE9c/DZch8PeHBa8iD9ry4e9V/ila
0fHIG9Gks17xRQKeAAU4Nv1QHYqoWQshl6l3jpkwaNgNdrglP6+1rR/+Us+o9oyy
d372clcsRdcCv0UpAu6rRc9K7CMcDaizZ2Rw0nP+gHuBo1SJNrUS9YVSg25qfCZ+
1PpZ68X/VRsSZW77XJG5VS9WnOQycRHGkHjaXP0DPEqB3Ru6it2XWyG8re7z3nCn
GBh/8fhz10+bCWqZA2bupmXKdjW8La1lWschOUjcqtJSdefd4hIsQY5flvfr74hV
OBZ+xIzvENtacHNpcaaW2O0e6kVEZ4FG7A5TlVef38vE7vFOS90f1MC76HYhcNfJ
BJjudrTFLWlv+rRxiJyIPkrSnCyFcqhkE5DPzdWh6hEYgK0N1cI/neG7OGDVx0P7
CTLnDlUrR34MhVqxdW9DzN9VPXldIJndgAwgaPHDodHm4F8kxmUN2PcMQ085il+T
c4P+/HWmZb/+kKLa5v+4xhplu6Ev482t4ZsswE+kmjr7rTHUdlcYS8gCXPS7hJpQ
FA8w2+ENlp4APUEHf0tfR4JdfixFnR3U3Irbhp2QalrxO8EMvvkTPW/eC6w8CNhk
+GxW0ZAzIgQ0OMeYkxfJjDrxq2/fJqrF7cnbk7UYTd5nlChLJPpf487uAK5EGKX1
qmF41DObZamgAfdBRh/BHgHXhUlz8vHRakZDQF6x9ehnOgjCJRirlDQT5qQwP1J1
YtmuIcJxJc+HsF5Th7ExXHNjGeY45NuBYRg4Ec6fN97UlgZqzGrsmLvHpuTfKrSF
erG+LARiF631VFyiFDHn6rk+i9fye7J8gRvoJXnWjcq0OKh4L04467NOJatlpyEu
yEGrOzPmbdLaEFiE+c2nFEoix5LS+V735nmGE4D2GahRr8eJwpST8Bo+LvRHhwvK
arDwnoaAfuJNaXILQEPBEIEVFgyc3bGkTB02jzczQU+nzgVUnBM08OgLDJcQSZei
ezwNm2atqB2kWbKE+cyJtmR2ogco7aMqW2nOZudkl6Z6Ur8S7FgkD+HJDXiU2wzm
ay3jaf8RPt2P6bIsOAau2Mrhtpt5XZKxwLkY5WL9HCb//7oOoCPoXrtt1qtBNz9U
KHHCr64eyxaKJ8VH0M2V5LyXJeey3rntO611wL5F/KwXF5+HgYbE+ssP9JiBk1MV
Wvyi23AfG4/U3bICIxW1Lu2VSTmKeUVvniriOpahy8BFF+2DM9u1NREb2bktdyZ9
TbSMIx0f9yrxrLaG1ImCI9vriBt9twq4PbDada+MbRG2O6SO2feLd9KdyshF9rYG
Cr4Za3gNOSFmYXOou0FAAdJj0G+MCDewvN0AXit31mKlfh7ZLF+ER944kGD+QdWx
3NUlWpUAzugL0hmtvOr9SBE/SsQw2njkfhu5Sh2/KBWYM5JaNUQqYmfJw60wV+Xw
fTxjT19DirXK7HEIxp6HrIZI1pXVB5CklVyJuarcRxMF8EK0LLl5LNv8E5bl3zuW
se8JvZYVVstDSGB2LgemXz5K69/d0VG3HKPgHuHRlDzTVp/yBQ9HzLscrW+B/1aL
uPgf0hxERVxCdj6JqWYUHtdGMRaksOymT5mZIh9abCeAefh8eaXyZiTNJ1QTZg7y
bdlGYb63eZUWuhFDCdRBM2xH744mBe2kCkveE9Ra8UBEMl6vkPMzaKumbu/2XglW
zQDdEo2hiYMqCd+i61ugcwZFHDz/eGIMXKQfpLSCTNLSKxNsMsPcduIWYlcLBaGM
Xr/xcvBDJaGny6t1au3qpjqDahNU4u/dSDszPxYvgXRKpFRCg95Ud7ARuydM9TrJ
25A8QJ8sGOF+7qniNhaBAE2RBAc1J3QlNsdgbTOA7GHzE66af1grSptj3Qdoifdd
Nfg6cga1pQI4DmZYHNsYgWKTm8ISALCVd68r10wYgvfC6OlAKiDrq+fUvczWUs7+
cOQIXQcVjxAPOy5X5TXxF/gZCf/SH3gvCySjVT6isf2kLX4YupChf7QYYDoNjDhG
d6Ut8o8OHg5NxIa8q510yQBa7yg7MIZBx9KwtIJBXcfcYQPMW4ulLQA3rPaoGHiT
eTWB+CuUfp+c+yNt5jePvkQI60pNVX24Vww/3y1qNUMCJyhpFxVOPMJv9Vg6+BYs
CG9cpEWpPBNWB3NuZjMLyYst+sv3YGJk0LTTgwVVl4jzjyeiCyjYtsKfLRA9AqMt
mkFj+6taCLYzYIH+NMykhTPok/0Q6x3BntCKLzTgPA8pNJ5NUyNyb7nVAZ5alvEh
7CoPikamQ2sqB6zTvWA+EZXX1XcYNNmfRaJYspZRNvuWlYoEwX63FLdJZR1MnnaB
eGP7Kspi8XYM8z8sn7rzG0C2hhUY1Ps5Ayc57ALZQAwN05Kh60uweCm7Ajg/5sF5
0hhDJ0dteXPwV/ULrCMLZ83cexsq9CWlblDmlhJsSMKqaLW1FoUqZ1aARdj9dLaV
OFzxhAPI08albE1QQGgNV9v1bSJ6zoIfEvU9ACrhPH0RSpUWr/+F8F4o+gOjG+rj
MhwalVBvGD09Z6iDf37T1jOmgfm7ogFFRAyos5Ue5uphsHxSoFIqIAPm8dLVW3jO
J/A4tDawdvBMDGzOsjquRaEERmwRSOZiQTMIxpkvIoBktXdIqHEd1fU8eOSMNChA
uRG9UuBKrL6F7XhKkqo6d7Mf+7Op6OQfuH2rZYI+p5kuC305AWKyVxKhlHmoAHVJ
WyeQfQwTVKeASxT8NPL180I9QDOngTleRum7jixciXbM95iulzmLFwwWh9wqK9WS
KnQPnpk/eDWphN9ktiQ+9Xz0C7N+V2UUVWLSa0DHC/043aQ5I7n6KBczJF/UT9rW
9/mhTde5D4Ze8qYiAQFAFDbg5pNFiwLdjwCoYwYixgXQeO1M7F9Ug7TXjdA1Ndbq
UuiUQZdSbfIhAoTLtUp/VAnwWWIkIHh5PVFmTVpe+MgmrQR5TPA4pZGp0tp0EEDV
ki4KVoDm1dl+ikeGb/QrtuxXLhNReEIfDZd28kKBPrOL166qeSmO0jm/0soAppZY
Uz/bbbGZlbIXNqxy0sgyH/rnuZWBDwf7Bt/zvyrmchZjHC24Kx64VPYzi0k7Eegv
eOqqVdmEXRsD9hwKekeX8dBeiam1xMMzjyLMmcks4naLfud2dkFvgbJiCJ2A2hKk
ewaB7x6YzyQe+YBOEl8QWhpVJmHHUWEJDpEAm19NqxYVySRW0srrjecVaiPdlrAn
gMGweaMbI7TCq98Zn1o5hy+f7d9VY2TazOrF+EkgtWjVjlYaF0XJNghn70BnXF9O
zOqhUvQTUQ/20OcjKhdgQ9/EF6Ioy1AHhJGOyRXSQ2goR5JYLTmVx4oDebNNqAJA
FZW6RPEXgZ938XLCE8Lgep4o30oyu9tWKXYTbvzlGN2X3MzVIg/iaCZNgtTaJmYK
DSenJbTyiQ8lJF1a4+5kQDUxeDS+Bx3J5Qo7r41970CUO2XazR9gWbjIGtRFCRP9
lhUGa8KOSc+5VBgLiakOrURyLXnGQyDEuWXbYxG82jmxwkGdQpYLrQUR0mQvHzZo
uOkDnDKKihHgiBVOTsCDd84hzbIUDNa0x4MN8kWLzgbankANgLzrUUG84lYJytzM
XyyYxNeSp5BGRPLRyllOFR1bw8kGPUCQWDpB83qpwl1uPNPGkyMAjz3o+g6ixuDi
InufD96mNFfYRaPCtDs2MEK1k5KWU9nLRF1a72wGz8ppqT9ABtbShsmV0xJbGQgp
uRf1bTNZTWKhp7yfQrLH49vexEKKK0pKHj0sn7AJsFsw11QXOJSZgY3X7kYg6txy
1x4WYaUfPntTeDIUocH2E4FYAL/NwejUvyxu/CIuRpK+tyjy2zzSwW4ufOCzNiuP
suUkpG7bsU4izNe4kE/7Cc0V27qTBMW65389VHbRVIRsn/TEQNgaKpfW1exhstFA
fMSB2mPrrG/GEAfswDpDdW6hL2xZfLhbZZfloI2kHxzfbPE683CRi2D09hMKy0PR
cR04ATCtW9GeXdEyTIyXdlbc8VdMQ5ae3GYzBvWWNaJ9noeUZVOQhS3b/fTJGxMy
OX1qtRIZX59ORY/z3CQSPNgvmpufR1jQKcRI36vqg+Yqv3km2q4AHF5cuDSEuemN
+yt1pyeH4b1YYZsrqKOGIpzow8P/jCICYbbTH2a6EC2Nt3CuqTEJ2x8DYzijn6X0
mjKC1nMY2UTNyIICfOtUSwkNipR8FlVDfMF3hfTarUKEijhMogIL+w67C8GWj2s7
JcKAvyf6r1MXO4H1ARd0+MMjw+ORDJSyqzQTHBdjS3wlJahfjhItZa37KaoVVm3K
pHlHy9tZv6v/tT7LrKOyZRaU5xz7SqjV2q5HVs/mR8e7haL/6NQ1WdHzVDkbQPD6
CGJDTz3W90DFoG6Hq26VTsJkuW7PP66V5JD/wIyCZtEBLq/PLtX8yiqiJ2d3P7+s
Hv8oqzBxi3dcRfhnEqQJZXoYTjJnk+9P79Ur2Uw3ufqECult+8MzPN5RhxgpnsUK
zGsbhV+2vZ2RVcaMivHxJryXLGK/GM8RRHNhvcvu67khoEdIilYfXr0KSVwYa8gw
e7wf3Flo/p8rf4pifIAZcRWufQbGcJ/5hc5BTpPeYH3+OfhZmXKkILe0slBO3Le2
3Cb9aLmpjr1RZWlN3i7zT2xGFu+SkP96LUEP8cvZVBDq2S3u56pB7I78ygTPwDh0
VFtSjNruKWtKy4DP7H18yHm91KKARAasOkmue5yVpGyo+d1jGRa7DtlmrOyrZzT4
J43ZTf8RQNwmzv4utWUX/yia+spk6jRrk1vvr4tB9jA/vlhzu2iByMujJKL3qrI2
OBbaBmDqg+UNKC/awSMq2npXS7+LFEqQpFl3zIp1xNdmkpm3hE+3H5ea/ovBfSA+
hcUEsf27N4bIGBCrKAI0XT0ksMoCizpLolLgKb6+4TVestPZlZH/R/n8y1B6/1UG
jss91hT7vgQaNiOzHw6ZqPdpCN9QYHqX3e5LgDAxlkhQi6igMmOpKaJF3Z2gqZ0G
+VrjCtIGzSgNLZkgvF+KTCug99b8oQveDZl3/IhtcVqkWF4zEYpmSyRE6ahGi7si
mAyGB/2XZIMZtzk5x3GdHzJBIc3s/a11Oa77Zsy31myBO1jld1k2FPlQadvgS+Of
nqv0VOwmKTsvsA912sD6yDCyqPRAcfjB9gQDvvsVE1oMVyNfwkVWXkowlsGKGlcV
qUcCwP5GuzYOmlv9GRgwEQZrLmCsdHElFfPndoUsXtdAICLiXaGTb1LH7mSgir/S
kdMMANdovEi3v8T4zYmjVfItc1nTQpjZ+K81KkQFmB3xYKq4joYKgyaj8eN3yXb9
qdXcfxIBlluaV4vuxZMrNR2YWxio3TQ7+SND4PrwYtTd3K6t2IakcvTdlBjTe9RG
lUG74qFkMEGFubQsmTRVAUZ0dm21d597GTm0n4l2QUDyuCiZ3eOiWIUZwBvSHy3A
SvLE/AkVfki7fCcq6cJBRrnS5DC9QeZM1ESo/KmJ1vuju1hRGP4VjbS98MGv9ncm
5uOtUv1OQXZGSwg+IjGA0ALr/3/Wsr/T4UFl7bGQ8Qb5c/XJXu8VmPvXRbuP8w8i
q5cQAcchbllTYj2ojtJNI+nLv65+R49gu4/SkOJlIfNQ2n0BtOftGQ6hpRUTWdVS
5ugGBVqO0cea9x39TDNEwBYF1tJO2FPo8VxiBlOiM4S7xahLpxXYD+sbwGqkWGEn
gVmbBD406RxHfH1cj8tXT49DITRFwtpwt7Z2c6AhYrlurx47balDgRwlfM2MNyls
J0+yqFRMyEv9nOe1xiK06qTGtvFYXAlIQBt7ucmcYggCylfNO8ZDyeJ+2WDJHUsK
6ye3DJWPzmU4suYLcuQ7esQ4w4RksalcuRrW94URyTBpgmheqYERBoUq1lt+5Q+O
abqk3uP7ROkOCFzttAyrDa7h///0Pvx9OWrA09VYywpaIRjaHFt+RZ7NF7TfP26H
LWpnFTKcDxpFyuvnnSpHvhaXxRy7ZxGNRWegg8leZNsu1qbIHTvq1pdYLVUN1a54
IO84FBsSAXPKmxAvLhBeag+XD70Nm6ZufuYHae2n3JkSh4ssPVmtEmpur4qjVTkD
RxHKvT+nrXIBwHduslJvG7uRfJ0LgfETCAHCo5iBFrIirD1w8C468hoYMhEo4o2/
CIYT/mJXAXoNf2lv5oo6kU4xvZ1Ng4L1dEKaL5JC5ZrrVLSmq+KXfE2nnF9BskGk
Js7S07LDG2RDaNYNQ2cp0ZdAmTReoxzJKZA/kdLfeMs4Etmw1r7j8LtVL2dsgWRe
Lbci19JLxf9foDFoeaF73aVqcZq+1VfObibYtHQg8j+XnrUvI1IcaLEnRI2wg3jh
9IdFPM7oBPjvdtUuLBMsN78CFDoGYtlj6aFTb1HfZZCSz2xaCT7GBlddpT+K4fXK
A4LPIp8VnrDD41ApOma/jaFwHN41W1kBDdsJQHoiqc4AmnOlh6JwEZ0pt9XUcFmV
RB2spBBfqk22EcI/sgl95SoE0joFIzKzNsmfQgnhm0W9L96NBin7OGxrl04lej0k
4rrGwwR2jJ8OxnG7ofsORN1sZFg46UC+/RkUseBI8Tt3+RZi1OeJn441sqMyy4Is
GNEBf3CHt5VAnEkRHXSGRTOTlODxXCFhmesVRgy3IacKAGwBF2LWnXTA4RS6Zqdx
S5Ur5PO1MWenpI8O/uHyeEsA3X7maIUdV+uQimtN7UOag0ujLqUI1NNWK/p6b0ek
pHsSitfvLxu+0tXYdLLA5aowoER4Lo0jGJGPgb5ZG/tn8nAg4+Ht2Sye/L2Dd8dm
uzVxtj734XDSu7SP03yGK62TD2oq71/4o/mZJ5klFx6BRoUV+kyJ+MXWWewQhzMo
qjMRATtiNtm+wB8Kd9V5oPuTIihyG1R2i1cHpNe+lYerRIJyw1x+oEKE+09ruPjN
PtIDdTOYcVTLZeVjPIaWem5bGbyBgFg6txqIIyTO2/NiaGyqiR+ibY4jcN4cAoQJ
38xK0ulgDc9RbqScPAHPSr+e3mjoPurPJs0udSCd9DMC55V7epgyrMNp0JPm4XXA
RaNIMVeJ3dzD45XHtIVpOol7etHz22lYScddRb8rg/siuramNfosZwuX7/4ULBQ2
Ph5Kw9R6BI6P0TyqMxXjQKrlXpDe+X828SULOWzDeUSz0TgLmB6SPVNkKCtE/CmZ
vGKvkgX2+RjrQEDNrgKpbZDBH0p81W8LTP3MyheeLbmH5DKcrj5pDVehrMwV6wLi
e0qfkvOEIRl1Ahu1QSv2DtMFJlIwYM70gOFEMuMsHe9BiGW1jBPTedhR3+O8om1R
ktXwaJ9dxYEVxbwtUDGKa0PPKSirMgpSkNih0Ft3W03sfAAq1Hc4o8Vq6Mkzu25H
Y6VLTSbRzxy39nu+UxNwPXVtTUtCj9lfK2dJx1mAN3Qv+3YUrekm+Nl/ZgvIYauC
Lnfzw6FP81EwrI4/XxCUKSJtnzwzJyay3n3dVfSLsPfLPKBrbV5kiBHdGe3Ad9PV
X+mcRgCrLhissB3+SWMmRLNdHvrOOaF+Vxn4OyFBJIgvtM6SmZspIt9HykFHzUC5
WZJ4C6TOeN33u0rdJIRLSc1NKLgBQs2XWnQvex0fYUnA/cR3nIVV35Afixk+FPs4
fHId3TJ0I5U2QqcSQRNgcQQEYEPtxG+14ho0/s9z+l4Qe7S0q56/OTpcXJWO8Mvu
UYHEPKQwHRXzXICcEBNl/tv2jcUyDNkfbxj9BNwYfafLGOVFb+gY5AK1cX9zaYoI
GvbZzUkHDIBv6C5VJne1qC9Hp+mLUTDCiIYyrjGPM/E/JvprnmqaNBn/hbXelc1I
UyDSrz+Yw6ACoxcLWtPlo9mMMXvotG808w6XumAHtpzWCo+E2qalmQOQDOsQaaBo
7qgsp1gb6o6UMA1OH7AlRx6S7KU21TO9glEeSarK5WLnPnaHbuxbLKifKwEy/suf
iUj2uSzJux5K2Hxgg5K/carh7TPZCG9agHfbcMSUcPnJWjr6AieD94Tuzc8LqnTy
VarTOFfgnQ32pfi7R0+Rsm7MK7wF/1E0RavLE0GPZ/RQS//Ilj/wNhSRv+kd6q7U
pOLxow7EGC5/vv1cDrkLUTcsYwDXr7cnYzNMQPYBjp/thGl2YtMezV/ZhByVmimw
fT4qSUpSTMJIf4W9AplRDOgUPSnbcob2f23g3uqgqxUdJPbjGUxhxA6feVyF0Ls9
vSzYvVam2rYRtdpHMy3/RQ8Gv8pkNwIiV6RxWrkJqqatKPSy6kIFoMO/NMfJVnVg
6V2Ooc1kw9Pudwy0UkVopcCAqKwyswDoJL1BVuuoDjXnXd2jf5LBwWy7tUYxx9GQ
G0ZaZYvSOXqIBdl0BjA6DqWxM0OouIo53FL1pB3ZihV6WAYOWQdZ5eDH2mfMSMd1
Q+SNK2BjQaxOmMbJZxbyN9Dj3ii0rFgCl+gw19ywRT8fi56cPuaaqG8SiSgGiEpG
aLPIonlRdKEpjZRDDNmxqFyj8VBdMVc6L7BBGDszN/qpSR7DYZO6tXDRDlzhlf93
uKLWLiU1S+MVMDM/lkRZi7B60Wiem0X9l01Jdv9r60F3Cc19KV9F7dmzSJzwKPmm
rl5tJVrjjgDdQ3UbtuVbSWxVDlrU9L3Fc/B20He55uk9y1vA3ijfgQ7gqX/37rDP
yQ88cm4wJn8206ryL6uAof7ztkB5yw7ZJ8KsCbNL39O8jSR5HyVwZLoBSfTuYT5r
8/YLgxnTF3bXVNhaXcC/WQwllqj8E7xhHRMU2GQtRo8r5BAvJpEWKVmGPUTgiVbX
sUoc+ll8upe82wwo2JH5kUVOFwsF5wkov0VK0yhcE4YHWyFQMYQecp4chp8fBe6a
tUwn42BDxECag/JjD/PgWpMnLEvqpNcLDgDFuxH45fT9CVMUUdl7zGJQNRA2RKyd
N6fF2mMAI0iBkfxR+KaBGooiB4siQdqlaUW5zTXjd/XEOOA+sBJtmka/55q9RmVs
PJgPDsoRbwxqkyfNI27ym7J4qaUFQmeEKAQsBEW1mfTu2mhfrsSTVIcTh55iVgoX
jFfkT1167V92fTH5tB4bTe1y7X2JsaRrtjJRuA5S0XZ0dMGouvKlZfQKldldOCkN
5tSJqpHLjo6EZiV4iD+9U5AerC3zQTrHV0iQEcUMGe1TCJBPe5i01+ujwFDc8z5d
51IQBUU/wtZP5VFrpu2qvpgyDNocVKHvJVBXypsKda1P9SKxm1bH94Fx/5si7AfZ
neSXw0JJKSfSnTJUfwfcuInHLcWgxdgaZ0vrzGnHfrvAYUNlWYx22jNoMFptr08f
495oyUCMLkrwcrP+RDPcu85XUFEOIW4MwpiW16eH3FSC1CufLa2xPm+ld4hesTaS
BpdwXsD2YWlDSTAtlniohLLtQKNEnORS98ngZL9Oaa48S/4Cu4Yr9BiGr2TOSXiS
g9b7vyjDXkdpshzvMwPdqD/jgTUXY4JcehYlBqgcjxwHhq7vAsdljaYEL4C7RZbO
qZd4+BPIMLBfxkIuf0HYtpx5gYEciPdgNcP5RQDpW7ADlu+gZp46+JEBuinzQbh9
mv+JcfMuxdoq6Ra37mCAJ9ErtHcOj7nMu7vOztL5kKTTeMjbrTBBNN+9lapQBOT7
6PFfYkuw4aSl4PN4HW+7ezyekhy1VDSgLq+US7RdOuSBJ8cZmfvP88C4RD4pWPPf
SKwLNkde7SPl9fHcONT14/UKhTVD8XUlSiLfrtkIs7leOpfJQ3XlWZCH79+3Bcut
3SpahhSEDW+VLDZBVTSZ++etfh6BUNmwKcVlnnqaNBXQ4cUS0LnldktCAYuQ9mdE
rRhLTYx2YYtX0db5SusC0qjhR0YFyuhgK3JAt6bMpHy11AzNWbzG4Fc2X3z+7v6p
SBPZ84lzDmnCMo502veMws443eqdcYSV2bTUF0HuhhShfGuU1iRvADYn8gnTYkWG
PyaRjB/qIwx0oA3Sd6vnTMBv0RsJ6KiVcIleGDmTyJsb9bekFhrYBQgNaRypWtjX
pKuJ10ER4Q6ntrAmvYA4KnOud0/2AounE0OgiLgDFUmRax5t4jJy5CY3FbOqtYPv
xtiITsjLMN0gVkqUrUD7otOUesdrcW9YuUxsQ8470sj2Wks6JLJX5JAaCbWWfus5
uCESAxlNf08zkM2Cj1t9cy8DvFL/KR2AJ4Ub1hbus93MtX5yMIbabhFY5HdYvORI
wxQQo09OeMqjYmBy/4OxonFpAS3DfRTD2e7zWB5dZEHmkENPKzOG4uLxEK4lKQy0
JavQXSmb5E2Opun2G4wueECDzvBpAx+lAxqiDs+N0F2B2Zo/t7QYHx2W6R+5FnOl
5PzWkTksGaRDmYiEVG5qSMvNys3bsu09+btGC3Wl5oRjYYwVAWUqMrzXj/434tg1
Te7pxyNlwHcOCUm/RZXHFTvLk9jpBOh8+XIdRrT7ak+9DiaJFv/8afUndh6FAEtf
JjCM+mqbD1zqPeAdk1SZxZ4YoFJ5lh8EM5T6Jlcu97Qp1IldOvTk79kx2I7NEuUq
7gEAH3fHDYIeokJ8PAsV3SxKsWhWhWyN36erkK/DipeTsxEwUvy1EsmC01cthAF6
yYz0G9mh65fAXL0I+xVzYCYJ5cHgdF9BJBk1QIrZGzgUh3rNUBz3hCfOhNV8BvAp
apCX97dihtCW3/C4cJWRkC1g8f44ZsjkLXOa9kAtJatdnX9bZB7Fj6vu86eLjFnD
iMzpA1FZiGVxO3YF8PvacfoLotEgyNuyavCW84a6DlRKILpspbDFNo0UkZYr35Lv
ogFOh34yahH4zixpXKI36yb2CSxqwmUBAzEdEDdlQ99JlQPu4qE8Llhpq669nX6I
4EJcJm56qTOV1OFy0wqvY6FB5ivAyA2/YqQfHqiOBAco/4hkcn+Bc2uvoH2Z8qSv
J3FVB2jxMwDx+s6ILmcMG5lBaBRa34SU+DIRCWUpq6Del1/7gpp0CjsMkr5MwOMZ
zXrJInCCLTWEh2niUDdGisG0Bf9mHyd8qUMP8nSMHuGywDkpXrDzeDghdx/7nhZr
Gv/ePjZUEkGXsr4/zjc9F8/Hmn8l/S6gTHNGfWlhPlR2JJQCYKCDzIFrD/o3o3x1
TgiaolfS78bZc1fg0dboVOy/3kR0k6QKCdJ1htW29MELpC0dRmfZcPWUUPNxswzR
ue1S2Ir3pPbrxyEXQQpKedlQYyNdjTyNakG6Ekax/WaFHsZx2ekXBIMEAqASM7tw
re9tKAQ+aIt/XALGfGWlpkC3PwH4PpJHBGbO1PlCmh1T9TujbOTksK1TIDDsGjuP
URqDQ2gg03b8Gg5EqnzbOfgF2Vh2pVHjQsiaL44gBcDsOAU4gbghAQfuzda6f47q
mxTzxudSxTXtMwMUQVDeDzk5KkWW8Q1/QTndYoE75rVW8lWket/6a1/UTegzN5Gu
wudvtCppig+zQe7oM4vVKrvy1yRrla6KophqkofX9KC0bLpgSU/hrvKpitkDuLDl
G2xo+0c9N2kVesxLy2KwvjfcJXbSeM89ormiTPUE7ypFQcVtTSzRvb0rgHzIAbdA
FgL15WRNBm/uRLsGqhCMOkKejRmpv2MUctz6pOgw9ytJQF/SO9e4CJzBLQhwqXss
NfMip8eY6m8GVMgmc36vmAk7qbe3+K9zEsURhaZk4nTeuQaGW28vNBF87nA2rKhH
UjXhBY4Cnty4GUU9UE/zixwwFG7X0WCzqn8oSkHAuSGJMtcPVrxP1CDuhHC8FxrJ
g3iBRzlYk94vkY6cLQxq86F09iWfSPW6+RgRig3/8l9JxOHsfka/QgSUOhtOG4tT
cfGzSduld69Z5AXTF3uPs74+UdHkvODte6Bx2DeNxr/tYr8UwAJaPtM7D4DSeBE2
Uku+kqWqaPuIm24+/BlOxt95ZjhKLpD7yRx0OIeQX3JC9SBibrd9ZhK2pFV8f4TP
QYzOwqnX61nW8DgJYRlbtc90cLx7nnQvGVHrUu/0D6RQ7Uiy+q24uOkPu9PU0CF9
a19lRqOXTUigPBE82RR0mwdtJpTf07n9XOe/YoYHt7zrxPHt6AJ0YpksmvlOtvoP
PEu1Bq7TPAl8XePl64np9w9Y3Zw1PE9RRdDM4t8576t3kUWG+qnBa3YY2Vde83ei
mY7Se7UTNvYX1rWr4MjE9LrwlAYUTSn1XU3PnXYFt0hhq5NuJz9PYZznDjrf2u1c
ZO3hMeNOaiuRsDwGMmGwFFDYMQRzJdoNEFf3n5LWU2j2CTmx5TYJgi2tu8n4cVPd
Thmy+PlqIXCb/emSUnoZc84J0YviiECvOXvjbgfI9+BFMhx97V08b7MgGBTrFbNC
OjC1L9WZy5epTdIIJTAgbM6Zn8rFK3E+Ut4AkX247KT2JmgjUIX/LUja6OCaZNn6
BJt4wo30BUrgShRnzliBGj7BWZmKn/TZc0q0LkinKbIpRcyBzcjPg35pUJhWkNS9
cELFQ+BYbXhThpy0xC+q8joUa7tL1k21AemUtWh+7sJCWibJPaH/NjSue1Fi5zQh
B2Xoinble5lTqqlHCEYsnRwfc10j+r24x5trCb4BX8+67xMYYSPONlQTT182On0x
sKjvxW/h1uIcNWDcv2fhNt/nGjvzRSydZ6mCu3/kYoxOvLA1c0uBGSf71qRwAakE
NIDGv0jTQTaWbzbNNKSZI6iWhnKrLja2EoW863pvFL5l/qgyf3+vKTEizrtC9glD
2CsfPkWpD5k1SObY6qW+PhLYyf7xL6WjsKn8mm+7T7EFcTD7WokSFU0513bCFyyj
NyjfNsyIz+Ieh2xgJ1DwRoxco8Nr+3qhbQkU2kzgos3hbV9AMaBNoN8cJdTctkmD
h7VFl4HEN5Gxb9Mw8SmqRFJtEFBtAQ0IeFQZcyoKqrqHhzSxaB1hRDZ9mSMdF/88
bT/Xm4ccp04cqXzrJhIagtPX31ZnsGgAeSFx2V0ywXLAXop3JyL99uVpHmDVatsL
YDvCS76ciiRiq/QoUkCy3wwPS+Tuf0GbfbCh8h5xsypAh7OmkLyTdr0+fI3UozWf
I8Cy8Fx7RMA65CQt9txaCPDFEwllsb8agDTUaE+PF3fNqyaHuD8CK9qGsZaU4f8p
fsCOv/czBRzcs7xTGqIR/v4xRlcAebv4dhAftsz9Y5NEXn6R6AJ+7X0jTpwoUEaa
XENGeShq8bZClkWH4LjyQZQlY+ao8BoDoH2Fwtdvvyr7zzm0+QESm8Dy62dTNlji
JIfvMGnNp10sQXo6yUnitZODHRFYDRpWWRqHNwdRhtoj+rpiT7yUYWujeUvE9+g3
KmYQm0DceoMPExW77mG7R8Qab3j+6qjn6groSO7hk682IE/isS4ChJJ44LigUTUU
XOvtL1vZlvVpJ2CO79DdZnQ/jjZeuwOL/asD1497XPSMZh+QZK3oq3n6TsURGSQM
+G6Jyio5ssP2w056qN5E43hLnSPtZvjcAlVZBTF7ZzgQE/QTdn9OtsxC36oRJCi9
tyO6iHURilvivY4OFZX/sLb33l3QOYx5PLPMQJQjaPagx9JduIFG2niDgCHXVwxX
XXutL1+p4g4Hvm9cHhgm97RidQD5N3tLyhmMEbwiKZH8sii+Im52bR0envfXuy22
6ES7Edlu2UfY6zgS1I7jAq6mpFfi7Gn7bHh5osQ5ZOKzsm95d1zgXe0gMUF3nq1O
QXbw6h0Yae+qtqyoBSAuwvDMZgtlQbCBT/gwG+3kc93wzjcg8aZuzv065wc/jNYt
eWXJrQhlib+ybXZIW+8smtH6LQJmcM0JT2oVdM8yHECzx33yLbftlpyq8aCNpUZj
EelQ4sLscf/lR5zV7k4uKCpxlSZFKvYM5JyGO8Ly/Ge3Urn+ekOd9iGS4+oAeGh3
4nno6CWKFTWLMJ9KBZAxyikh5VZEUsauBEcSMoj17eraLm2g5KykgqqLX6o8G78Q
q5zp6B09byCBpuF0KX9mDBxHqPjraJNF3JrZHuvCGQXV04OEj+GfqAX4+6Rs0aka
q7GBNUCmDfdyONRMHFxGkXZPd/NaBA9qBQgLiSmio4RTXbSkaBWlXBGUMFjPA2q+
TRabpnSyldNrBwJbV2rGyIwMiS/+Ing+IgIvutSkJC0bV7und/iMbuHpdfzrH5S7
32f0KEKbX/eOekeJGF7GpPwRrN53r2YHM6pRH2g1rgufmcOtUSZFWR9nGsrZ7aLW
DN9HfiS93uzzOWwmneRneaWRRtFWje7LqfZjy2ob3RC3pWVPLtdrHz8n2WOB8XNu
bZr0lliK3uEVyDfLErZVt52E1CO5Z8mtImQkrWtDTRzCn3uCxO+npvdi15W142/J
jyLFhBVUymcfAmeAEIRheSnxG1KhH9yrCmGi8hnEgA+Vku3jnmBX/XzRvcW/qjPp
5kc7dTJ2Ba8nO9q1A10BbMl3A++KfGQ7MCQzRVzFq6JJtZmSjQXUFGt1H/SLb4Ni
2D7rBQ1rrDSrolqPnYxIbu6n+foj1pkCgg9UhjSG8y45nVyvwTAN9U7H2TjuTcFt
PuYNcra5VgpjB8IOMRrA1L8ZEhpM1YQtTF8herSxLAZxlUd2c70QfRqTfGXuYqgE
mrRBHfu5QOJYG2BtcmZTOIwFm4WVYxLbQHMikAi5baZInSyU8XHfxWr46Qbg7Fvo
RY5tXKmL6HXUEkWcgpxbxcYQIzfooWsQ5mv0Pt1/MUnf6plzpq+GYnVsU5Gg0ioF
QVVozNkLlCE5eJrqFsWHOFEyLSjzKc9nE8tzBner65S81S7VFWHvrIbXlVQN6K6L
0AjEsDLu9py6czq/q6EusNFSbwgK6oQCjUgOp0RXEhqfnkskY2S1xFBS0rxzNI12
zzvUnJtqAfZsiyxRdTK5Z88ps4FBchZkWz+oT95ozpLkzDPKKHmPoX34hD6UYpt+
7ckQSMq4EAc1nuqivDtL9n50M+MqV0taqL8wJylaENMyG5ZwMZbd89w7U5+1qmRN
S4f283u8P45WM434P1qcgvDI+Em0KDMe3hevsTexEbnATbQ8So/vMAOhHXU0hP/n
V869hC/oC5pSddpy9j5Re/VRS7T5fpL9PFLEFmlZnbv0IVq7uLaJ6h3LJSSWzENM
i6RO2uNHxGi3lJtAG1W2y86ao+0WqG3et2/QCBhURpAQ/qgD9CAZzkQMN2cZjkmk
0kdA88UwG3Tj7Bi42B1pX/Ijffm2gn/7PELJVlKfmRDwunc0J60tWaUBP3Lti2Wi
d30aYnuHR2zSojgAQ/AVh+7f4w5s57V3HV8ONdgPDrcy3eoELlJfwXaHgehfskKP
52QisZk0tB/5axpSC4Spfr918zR7qA4pwMUFem0e5sxfyG6O4PoRU5go9J1dZbPk
Cf6LFNIe+kQvB0HZ+d+Wc4ci/ACg6G/GIolK6Z6EOYqIzuvTgxDg6yrlovfEV2Ux
AABmlUp03Eqi3m8k7neDp9slx4ETbuDKQHqCZxzNHYYA1GG7e2q/9kAMEdWZpRlT
WAec4zAg4/TJs6yHIFsvuBnNN541CXcH5PXAqqxWSa0Y0OxXj4Z0x+bNjopSI+PH
N/cJZ50IkUUJmY20BP9Vnfix71fl3acaqhGTtiwE6WQTwR5wF60W9OMdYozWnjDb
TFoK+dgIrSzZZCsDF41FtNzb1ALJMOK3gdAgOOEb4xPQ3ZJNuJ+uPa7Q0zxrthrh
zMqlSJL8iAKJJTclu7Rk/sMsP6mppk7Ynnj6rW5zPuc+VuAd0JoU78cU7fma1PFB
TXKWAXUBmho+OOUSj6MQ8zhxFVTTQQWh7169FJ7yKnJ3bMM0E8+15UsWCF0AS7LQ
fRGsdWTxC0y6s+mBMzVQgxMtxHevc596wCaOK2PRoYT3Zcuwqver5svUgR6Kwix2
ixYX62bs5xUWjXkL6YYmcCy+3Kp7Bi4AgerGEs4SUtYQPehYw6CnVskouJMzc6uS
lmR/1i7pq26hYkiMYszfoN3pez2I3TmWinv9uLBgxTEQ91g5fqZL1mmkB6qRaoWR
foXgJ1DKzNPSJbMpgRJ+m2wCPI1ESwu2/OKxjlaBAa5rgJB4u41v+P4xMjBExGXa
E+mnoZ8D926AyC65YND7+DZuZ+jpVwUUi+V5slPBhQJxw7TYMn84Fq7Kyj56mdm5
PP8l5prS99JTq29zEUBIQuQbJdMdqDbCFOnKDh4BQvH1H1zIE9nGTvQLuICRR4Sg
UgTnew6s/g6Jb4UkDCgHQBYp9adFFJ7v/fYLOjNyqgeg42tkIcsFOViFiurKPnsJ
LQ5V7q2v7sQQ2EBUpGmqHBMsgNKjZM48h0KbXKh3sj5pPKlzIMP4UwrZoaZfC+sG
017CokMUhfr0fDQXP0HD63Djgi7hY3YDHO0YhKY3eQp8aUIM4i+06ztGUx2YRyL9
Q7FHms/tgfzq96Z6YSUdvgPJl22ch64DslsAOmAWw8EvAqLyg594l1q32BCLZ+/R
doZJUmOBrfghdNPerc6lU1Xkatly3Oz3/mdO42DHqsR+gRNqP2mbxuQtTLf7nnsp
uf1pRFPDI3RoYH8kBEQz41MliIx5412UIWfiGE2e2an+6/99F7HxQ/6W9ZV1MX+g
01L76I/Q7KIto7vFzHK8fZ6NL0IxLFE/srxHmacZ0Ouf4E1nN/t7GZChtnyvIDU2
1Y25pb+DeH9y6q4r4XR6HWPh2MZVtwsbJzcKcCuaI0V1CyreR7g0Od7R/dPjdE8y
Qytg5DnB11+jJllx+MkO6+RDRIRCUlZNBvtvwdjakVlS5/HxjXfi5V/55AP9Mp4C
yDD3zJJlXj62jSg4xffQV2TyZJgFcXcOfwDA5zqB4WiiKL0LzfsI5JgJMIY9mQtw
28fYLMaDnFYE5BYYBSwBe3vVT4PP4DkJ9IPceEvMLA2ZJuJPHyCuNdADvaNAc3rR
RJx6zYjrwCtTS1BvaNQaKXDBZDMonvccteVscOoXrZcicuFGzgxKN5b/A+Q6rb5F
UY8aBawk4DCLsxf5B/zEJ3A4sAuGMlKNIJhcQiBea1L1beZniExrBzOut3DBVVS8
ULNVZuJ6yZPv/dAgYO4L17FuvGdeL8/VqKD84dRyRsYY4tmFIEjswTlD7O+XGYl8
S6LDT6p3VzgG3O28P3x3q/TNW2mRuD69IZCk7mzCQDOsRyD5Ox0ipGzgvF2kbcTY
3kjwRQTdxqfRoci6w7sdWzt4IrAA1Z2pIT8S3xN5xeL2XxChrdCYyQkTbDHjZKDI
00cIUhe/dgeNmAmelefm1v8b7kjMJQWhx8dWeWWDesby4o5JsmMLDL9YfBIv6ty6
MJhwjnACeCh/AqIXnAFjDQAQ+xsDYmRYxHhVqFBM88a5r4NRwptTzRBBaP5g0WSD
dZJT3MTUGwxI7VK/a/fu9ppw/83qKpHpq6dOsw0TK1O/pcdVDIH35xQBr2K6yN3q
VCx8EIGesYtrAWQVOne8C3tEq4hnd82SdoOqW2lg0QCw1rWV0PQloUCqMK/EX/Nv
wvF+h2wYEaGJhl9iaVxs1TOP0ACzSMOUiISmaF7CJkXPC0yAHeed8+H47tEprjme
9pEXI2JC8F237A0SqhBvczcAwiSY4UGyVEvfur1gKHfkPuq2l4/iSLbjZtpkNVN7
pO8BL8BSnjAISz/yfjsA9UVbZe/S+MsOEMKK5gjp+V21zfnL3r5sLVYOsx81hbUG
hweHVcQOBvm1Tz191Lbw4a9jMd9eHdaZcu2FC8ITw4b7CKdX3wx3J27X0oy3EoUo
MpopZr87DIa8NqVO6Ay39+t+SsGAyA+fDFd2bBaPzy+yA7CnPmNEwPybItir4oKf
l4wbIH0e4G4CaZAV2HYqHZZbfahi0kcLPHjAXUi3e48qW8yhEWmUdaelxAK0hEQQ
5VOvfoccdKn2hZJU2uQwg27591fCnrv03SGueYz/SgTa02DChJIwj8f+y0Q3jiln
RTDcO6uRmNVCHlJLQhsKouImVbNKrp62ga9Zn/jYyDCU1I+dFe3NbfH7t8EqNuEd
HyTBAob9BLB4y1VJe4r3HoDKjXW0hZUadADewXYQKG4OVSBjrMGgD6rfMBpOeQkN
uZL1aVZWebGEdMKbwDwuqo5wuTnraG8MiVng3rIhQBqlT0TT9yf8z3rjHu6gbblE
l5UrETkhNsFNDikPGRJrkoWfyqCxwZ/HsfO1Th46hEzFFFImzHAsdw4qF5O8Z+BV
Y4YI9JSKu0y22iCm9RZs+bwnVjkxp2m+gHea+iRx6wuM8KMcEhSPLAWUT8pPjBqD
o5oYbgt3M8koMJ0xsukYe6QvyuLUvdc4XqGAOTlzifEaGZPY2wK3EZ7UubajVCwi
9tRLffc7W7WAW1tdkQfhGRD91DhIg0y39tJST9LOQIY/YtjHw2VtXO19s3rnoi+0
2QMcIp7ByFh8yQ5eR5Nt//QpDWHyAPSdyab5uYe5n/2Ng6oa56K5ImKjpMjNK7h8
0FQW9sIZVJ2tYE2gcVUybr576roE6a6qrP7DU1TUBc7ebD6PJyHdWEh0DKuWUc/D
NcmKPsld2nbjqvgdSZeSkxH+JuMscLLT849EdlYQrfhGvFUF1s4BBI3RIspIc9gD
ewP/dKT/fd7RitzLuQ6/MCbYBhuqwAt3d5dA7NrujJ7aLXouUFFSdQyI78ntahMf
m1XVla0l4vY3Q487KT5HvpuT9fCFlX1fGz4pj0r0NyIkvR22LZ54jzm/BwK10Zd/
qv7QzWiSQrRzDTRahxifLzx+JxRWNpsSEst66dmWnAXaZ2nD0t9WBKDxvaMzEqdj
LpU+WiFAJ/WdHM3UAZDmaEiZz6KSKL0tC++2rHr1ijZpgHAXBl4DMQvH8dXqZcD6
UslWEOOAj2RpK8V3J/2ojVxWd2Wd9dQ2PBzLOgbix3Bw2oMPCL+9T1OsmWvqgISI
j/x6r2pO7UVTrIas4zzCWTZJCjBADKFF4E15/dZInIR6cJeB2kEqviWxaqMuek7z
DrFhpswvEiLFxbhXeyjNTy9F7yN9CXAiZ1wmm1zCnDZl8HQWESSHIjejRhsC4HHJ
Syuj25U+AYQrP+ZviF7lG30YLiCcBNwhTOlfTVMBWu3PADJzIo+x+i4pt3mc0+PY
yO8vHeEVnUp8+6D33PuNTHmRMFd3+RrdJyMnG3Jl2uxKqVvHaDQ9LMNcVDAInK9g
Kupzez2Jly9Yhn6/WmxtmnOEwl3+AO2s9hO+IhxL0VtjLeSWHG9wTUZQZxl530x0
FDVco4zzqP9dmu+s+x8eb6yssqZQD9erbt5JjNxIu/rYAOMfw112jqpQ1qiM4RMU
syB8rPEFZ5fy++HRUG6zAEjnDtAGW2sKAOf5FBBGocg31UqZYwC3sf5cW2xM2ZY9
vt+7YVdh1vSxJ+Oukm86lhkBQ9prVUoGJTdy15tQYC4UcvkThbEPVIOFzuODahPj
gbBNHpdLZN/fuyuYGdo/jguchKbyzzbuYWmUg4tbwRtkTR5QL6ObDGlOrd6qvyt8
7xcpKWwE4oTbmnkmujICkwIm8xoY/VhPlwLNaTesTzU7SUg+suXRp9ESwTXlX4i0
wZ86kms4Xrtq1eHj8IGiFKdNlOGanpjS+yiXefGUARpP8WKEV4KZZzZ+gO5KE+oc
A30cBgDIlGFq9Q6I+HbEukOUMC4VhT57InfMxz2kGqn9dVXFExMv1kC/iDC0GfhS
Kdjw/CyLfNz5PgdbMkhKt4iXYjv993+pu/VqJpR5jGSoaZVW3xD3v80nl4d6DvKQ
TQC9QcxLXq/4IOaEZJ4c4jleeMU/WOcQOkvjMftap+cy36h53tIkpKUPkxrH8QAP
wOjiOSJ0TY0giOXlaXLdRvv66VkQtnXhFcx0Tlg8PjwsnaM4VRbhIZT1YWBuXHNX
L8Z/ls35QcHu5QeuK02zsVzb8lur2ZluqzyoJkQfdpIUDc0dZN1EjRdKrpisZCNJ
jrc22OdJPW8zYeHg5aJ76RfvRIau4GS8tKjgmenl5M6DdNdMNaTlyV1m8zymfN3I
sGzeKRdCQoaScTS78Jw6ggfN/DdalWo/3mKR0fQzsWGQNAQsEo6G1fWwxkAzML01
17zKxQIWd8NrhptaGjrG8MMmh6NWMvHKbo6wiG5dyy7bOwVnU2Q4KGQGhGUD71Z0
cUya1dz4BjtoQ8PJtNtamIiyNQQd8EZFNsPRS2p2zcdGl0s+Quxxhz4XAXNbXQtW
niiQTEZZAXNBb/fvW+PU2h/NtHKKGT4qMee8lAb+8RQREzuKthDT6AE9sAP7OM3U
vUQuIFAcVad8PJzwA3UVHXNQPLLi5T0QZ8kgfB0DGzaxDo0D8f50KEBl/G6Yi9HX
7c33Bafa9tNUXhAloevM7BEeiK013PmVfBdj8FQrrFXEIPDxgAafLf9/VOy1wFNe
h+faq+W5zBm6ZtzhxScw5A8uf6ADZgXiz9JuHYJrQ4WdyHmeHt+fTLNm0LhLOrtB
QqXfLN6oB6JBJggWHYpTtoqkZNHyqMpjcs7NhM5z5Izt58AoGez4sYuFvik2iAWK
UrqnvX+UKoGEm/Nv+KCQkq3zYoIc/kAq2DoypEiUknwruhljVVcTwe2U7Ye8sSYt
M9z/26ZWVIwUFiOFzDGbsDWk4blD02aThPfWIFYudX3bCRQZrqfTAZl34HuIYIJX
inXSlvu6o2IH27OC5Xb1yrlPaLqupdqoVk2144zxlHsuzn2B5eYBuvukADTCxB4G
48fuZZAys7XOHOGMHOW38Js36kV+b2Yyv/fMY15PUQxQs6t//M9KjiWk6c8zQX3H
54xRGpJd97erJvcEcyH4PxDpqfXFAbhzaplY/ygydkXAuYcg5ra9+/DXjGWQGZMS
ePksPPk/pmaCmzu0qaxgPfJ8QGPDvg/9WQU1BDYkX69M0ppnsFXJ1BU0MTLRe2Ji
WZjXR9LbILaSS1Wl7A7DcjFHtZXZs2t5y+3so2NbPn9XALhmkrAXYkz34wkMmGjw
ei9+Ku3AkQAdbylnhtS5zwp+FbTY+YcqpBkWdrIFaIDWwJ8pQP32QvxQH1BkXeRk
3W7V/7742xcwsAqTNJRJ5T9Z4lEvqPlibiqeyOHFjpU4UzRoD57Scmzg7INpiaxC
sFOaswQn0VjdIXrv1mDH5Yb6CQ46kl8hE8zMixoTEZ4ezaJ8KlXX0VktO84E2Cci
B8m6j4DV1Kp1iL5OEB/wBtnvfvm//orLJNGR8ZppmMU8Q6SsrNWHSsupbSMz76Cp
v9xBkFbfDHFohM6b2o4Nb6TSQ0OymUg2T7ibn57E+RBk2DOqJVwCYJvmZyVLWAH/
jfWGZFoNjOUHSZO3pK+whhohqGOiEr9NyNE2friAK3PTAEvcu6Zk74Rm9juMzq0n
rxoW+dnihNVp9Gz0ZPV48R7gV6Ng+CONRbk2cK+JBZQQOyuVzLh7xxadFizw2M53
xdBGY6+vzJQEcVi3O1PNrst7mt9WvjnQlhjVQRXoOJDRKpki9sYAs3wzz+ISzDtG
ax8Oe7nRWrJt5RZRPXDl+fjufkwwsNfpDn0jcICsle3bg8aLGrCuSZS7v6s/zGbt
AEHlSyItclZylrrMItEzZy+TKCTitwL34rBWTLSemItno4QvdZyO0jSje7l8AO1X
pJR3iI0BqJM002YaPKF2UhZDzejK1rFvJXneoxFo++G0BeUsVgOtXGEitk28teIZ
lUwy8rrgtTP3xCqou5ga6lY4ekL4foaHy+gl4q8YGaPzsUHPsKm1usiO2GizF1UB
gqA8E0rOiyMUIx426jiCsokMLONsrbQlvfU9u6cbzXgSu3volq5pB2kWasPRNGMI
2t4N08T12ae8XkJluJje03WoqqFfeHZvG0erPUDWe8BDLgJO4DrhKw6f1LJfZrkG
UtwPZe9uc+QMSB2zyZ/dzmNWRyKGSnIUn4EFKMEq3GOA2IRvJ7Il1oYY/gNjxBAF
Do01lamlfW2hJHX/wBKQbgOW3KgKA986YdduN8kJu0oPGSshFol6J3InGtQxXhsa
LV8Wxqov+lB3TEbVgtrXbAYGAVoRLWcq4nr6KJHDTaW08BW6KahQWLfsKkhKwyDU
UXg6FjRDIR77LV3TJRqqdwf9CFZbvFKCySb4xXQf7+J/LRru0qxhEHVVRQ72vmjs
x22CMFnxIiEn7oCBbGxdI9Chy+iD+S2A3aRFrbcNZ/ziLvqiDtFGoqSK+kjjsRtj
yCwbqVToiYEx+Hxb3WKclsdZI689j7u5v/hQs2wNFsdUl1f9LWBoXTHcD5hgo1kc
AWeEt+7rI8+24sjIdqbZjCeGGzSuXbmnMHuvx1nLQc6Bd8tV9LzYwj4gBqkxTKh1
xaHbLtQVwuTCYkslh8Fv3R15mC1h6PKdDfry6BB26aEH2WdkVQ4freqnDWOMEfMO
WXI6zn82WjZNB5qjD5TSKRKTIOtaAYEvfOlSIZ3ddwR0Z4lavhjZBaeeUinM4/Cu
4HZUfoV+sNkTTYtNnFG36aG6sxpoYXi0NTaaTDvNEEo6QmibasZqw1a3bP4QSeWu
XDWr6G53068cJ7oDeF9bKUEnXnrpWe79ooldKUq32kXfkq0RYky2YWwwVOVrv6hm
kua9lrUgpZ6Ckby/fU0XJDbjULSH3RUSGO3IDv9MQbA48SfLZYC2NlExucfrCWi3
H7Vi1xA/Of2EgQobH+G8TlCfOhuqfdKjTJs59Lbv43Oll+jYoHXpBTE7mK2V0qk0
6NkjPg/6SJZX3BJRDxZxmsHfZHPpUoVZcMmXIFBbEr6vrjGM/CWVbXf9HQvljBVX
wWa3sdYg945h0V5GAZDtzdAJvZes3wkFZxMWym99yAJjnsmvrXsq6RiK3rkPeRyE
WdrgTBPPdGf64Ok4Cw8V+U6+66KU/29r5lL20w2dBc5VT9PbI3RUNWiIshuNAlgg
uSi9gg5Kpzmv4GS3s1nB+WNJBRXqEeQSdc5OuD+JqvBaHmq4QC/nQFgy6n8hLXee
qZhdwOJkM08xxUrHlGJyOdWMRFqPATET6f5tPXFoDA2Phzjpk6a5GLY2spoI1MbM
uSID45puSdB4IyDrY8h77mXRdO4absvq3WQfj5DUdrUwPhXEsT5OUxvU09aayERz
pSW4vO/LlEOl/DWMf80tVsJESBWzNy63n6/Zd084YL2nq33xn4G2BVDvTMqtWpGo
IuqMBNCfb0f9LjJAFVZ8xeXysi88ZRviesYQRWJhfMs2hkWxdVZvu7PLxzVe3oGW
TRS30XcyB8c1GhYNUgkWWiApv6TwpazL34hVJd5EzDlMAd7aTcoWWRTuCIwPjoN9
SyKiFWmMjB8+TYnNsNdyyoDV81mZJLukXcVOBu2SNboYM0B/Je9lBLQhwmYJmBlu
XYRrlWoyK5YkQJ+4Wb7z+pc/XGMwXDAd37EbncT0fPPcahMvKpQzbpcDQQKZd3O3
LbLTZZ2zx44ww9F9zgAODAbQHSeltmcvhtUUBJXxoBFI72RVeexn8icLfpISn1YO
xAoxSlsSCvZWwpSy+9LNlh84jCWNVHyPikfXO3l8aK5kxLhIXU/Z9FKIHMH6o0Jq
oTGOjO+N5Xs4fIqI0fxz2/UEFvicNS3SSAbzUOl6lhz9F7+kM9AkWSV5R5oihY11
LwQp7JkQd9tRhY5OH/RzkVO+KvYqziU29Nmd84ARLf+a3vIYD2rn5POxG9HQLu0G
RpY5oOM+YHP0xbULKEZMiqE0DugfmSFuPwyGrZt+Bix4sOftF0eiuNMTwYhvmSVR
Q4DqK705lmkDg8tPIWCbDaaKlJomNSdiP4/AUjIIMkqPWIbbQWO8Rm78pSsT5miv
sJ9mx5orvssLfvz0/I9s+hN9rQUFY+CyMnLbyfkJwws3TXVFv7UMLv9w5VGhz0Hj
QFRY8goDzBWdxL5Pe21s/SFZFgRF8tu+VKmf6fUUqj56S6rms4CvFNwlaabxBpe5
w9Ye4LQ2R63Sc027kPRW4EPuQ/XXvpObXbmCERYZz4Sdtku96zbi70lLc7oghqCe
SSwDdp5lCt8PSxC/GTD2KbMwYTlbgcxEnCpMRfcvx+k2qu+bHOL0n6+oU8ruMs/W
LCcqteCyxLBIraUPNmWUonICRNbgUMJ3QchWKPqq1jiubvHpubxxqnUPs38MqWYH
AoWIm6c39u07usMicm6yyo1NdMA1N/Favlj+sJzt6eGJUvQXTLxGkj9fhqMOns2e
sTkCMS50ncsBN7A6OlDX8FVFyYRSHD21fRjvqQCU9vRaQVxcxNI1h6Q3c7uoWEKM
GmkQ2oFwlLwmGstXxIDTC5Hs3HNXY0k73vDXKZzpMyU2dePBS6ssfHQFXALRUBjr
Wd4CXWBo9hPufpEcQ0+I8FN1xvO5aIoQAPOIPFdTOJcdUjNz5xRecy2YQlC9D4yE
cdTWWgzsAHOPtyAlyfUnBZUIxNuKzpPfFx0ngZYta9NYni1tXfe4k9WvSUnMctQH
ezM4E33IUxE/6UhrjGSF32wBRObhRxghmD+5VVAK0FhMc+c+omqXXTC/HXbv0T2F
c8PuBHPrF6e8TRfttMgtnXnYv/k9Pj7ZmO3+1dymiq+yhsIFS757cmGEywSH/1RT
GU0KUQVtik+QmwAz4SMhkHP2aWD0ZWZfWjXMGSHdP7SxedAAc9E8ltPBQQeS6Q3Y
sELyuzFNLyKGS90F0lY+I1TYvzSzhwfW3K8hKiEnbjeV19hI55+K4RbXh/lNSl9E
6h53GNXc72Omhjw818OTgBFheyXe+pmU6TjkWndNnugH76+3NDKRh49hmVxoLeLq
9hdWBDqEHWKN1VjJrwHU1OkK0ZI/WT1EaOfGZ5xXpVtCVntzvNteaaAyMtCdmKz2
AXWDWMWPCuOuW/Doc1OSEMjiutktYVbK7uiF2uCBVOTnkzaVpmV89/gJ/sBXbym1
q3mwwyBKZgS7mFfyXt9GBraT/ZpRJdEZIYy6F1yvCg4XOhbhhSUiXzPK8BXXJmQU
qOktkXc3HRlURdAsIq098WUr4rjzdJGX9KIiIslAgJ6ILTIna8u9VGbYw6cnowYU
IxFO61hUn0TaU3AAW51znAzCZcwhLCLBCC/G+FJpyO5WgSYH7G+03BJwt3hnwMMQ
LlGo6L7jeB/h1XoNhCtE8UCy4SviqOjFjNcX5RmVk63fn6fd8XrDa0s3JWtHY0VD
0sM7Py3JNec1j/Hj1UGGHGO1cVMvAmumFRFKo1sHl7b6UviUw5nVSUc8Mar+OmOK
+3KKdNya/ELLcKrmPFve/c18Mm6FtJWJ5JrPh3yPqAB8MWNKvTliDCO1ePfGzwgl
d285GvKx1AbygR7pbYe4vEry8AoIXCTaSR3yUaw8FNwK306v9c6/7gw/Fgzx5uQW
EbN7u0VDbyPufjSqokZQfT+AnASXYa2WDiuDg2vt4fDZvWLTd/ccsqEYnZGXXbK1
A2xkRp4PwFtEeU2aB/4NeKue2AaqTJ9WwwpSpnlVfEN7A/Zwxo8r2anHe5TxrUCt
3GCSLFKkk/kn3bNykuYaF9atCSNxe9pl1ZUmv/BFJbcDpFC6jGYmhBHDKsK6U/QM
5/RqMLwl4chvFzf7DtkRgsg1FI0hJtrzcwJox/hF4HS0+tt2Q2TF1l7jAWdCUv5F
Weqs/MrrCQP+dPcTKMDHkgkS1x7n+SaGbHA1dSa/mV/n6INaM+CmADHwdId0xmk0
y5hobMuBIL+gT307HFrfIL4YNg20KKI1JYFFzu+Z2Ff3JRHAVr7pTiXPdoowBWac
PUhOGrSiQyw4fIQW4sT6nMPeb09ve5R5WF4Pf5bOMwJSKpermK0Hf/U1vBwBSkEE
zmsUUnpxPCgQM0BCLP7KtwG2G3WC0ooLJlGpcP/ctI2B7HedTRH+ciJwWE2Jnx8i
9p7laUcVfqa/ql0l6vlf9rXfjrwLvHmDf4p3p71KoTvldgs2UxjCkzOvz05vus8i
4hMv86ZDMaVcswc8QnzYZnmwhBPUuGfMRvGUWLTq/+elkJnqxf41LuW5oLvDEumj
A+3rABmbMUMB12zx1/5DFVDMFfeFAlnlqzURIzIQ9qd8li7VO5+8UwA7iUYnmMe2
sDJpEI24rO0AH2gxCspzTx7hRMaXh/3NY3G5q7zg3Z8aGXDAJcQFiNVP4eGDAm7a
K7S/E3K8dV951GAlD3uU3hfvZGz0bNoeDELlpfPMeZkryyyymGxTb4qKS/GyH2Ln
2hKr1mqmhIg5/ChqfbJLfZHjWIQu8ggL2nL7eBwG9MsSKD6/z9GGgCulS5KK8OIF
7qMtmSTGjbZJAjktl2h+deJKcOaYQ8V12CzJBFhfYWs+QNn9E4C56xdhvg5YPT7e
yMUxh1jB7VQDXLSBzT4hTCqTKG7SF0STiQxj3yHOkcf7fdsG5EzKPNTFbiTUDIC6
68OiAGJ0IKHI+Av8z0a7njZqRoOqWLvvTfbhvQuLNsfZjBe/b66bSVaKlT+CiYq2
GBk0CunGdBS13AI+4EXJPJ1N3aF8UQHrvNzHry7CmQtkDa+6OnUlnnqY5VHVPUsJ
gjJnpD1cGsbvSH0bfwFOizOm7BiWFCWy7RU5RzMl09XrGkmeDXd+E+WygKCo13uk
7CeuJkTpfY1pss3cjxYJQJu/dqlLK/gIMb0RKpesa4yNHqQzrHGR5c149n3bsrpc
DJE5fRHPuptthNQukGFSXpCOKX5293pFDb/Y3t2aNvbQ5gEywC45Pg/b4Ua/bZ4m
GU5OXTF+h7KNLsqSQM02gjpR99D2OTdcyPTFGUPq/QBw1V9m6eD/Yjvp8VJBmHP4
n7P9GfDZpcWSXYOEwhSQ4lmUNQJAGxmOeyvPvYt+qXCCDtMdMHCbDqqHfnSgM5Of
E/dK3L1fW03C+5s3cycWtymdCC/pndBC9ORdBl13y0NCl8DEBBha9NkX7zFKF0UZ
xHaFIpOQfPN9DvUGnkx8KuOBV5FbD+uM7QkrSDvgeP0ltbzwONf6zN4norz6qsZk
GA2ncWbcouAdWcTwqlYVPQ4W+zuC1+R8NCA2YG4mBCWsJXXAX9YCdbRGVqxloKcc
M3IDfN4j5XYAGCH2CoKCequ90AdrtQl4YdZJD4qukcjfYlWSR4H+q8G8jWqKKUJf
8pts+VgZ5IOUnZdvMfCkg1BF7JbqPJTjmFQutZSZYvQ9exm8/oTN770EZFFrm9hp
JpYgQuTpVGVz2MzwtDhwZsOnV2y4SY7rG2I1UGKLUJ/3GV3r1idaa62JE1KxfYdM
9dxX9u0G1BFA2PiuVz4EFqge5oGxfGgaege2R7ULrdTLywqE8ahIYGt7/t3y8SLX
yE/2A71G5dMM6DCG1WP4vZpoeuo53brIco3gIGCt4Zie+pU75UyVAMRr9a8qoHHZ
1jp9JJ9nXNhzDiu2jTbeC7mMsLnHJNqdc2+RuTAhWezIY+55ISU9uWeqjqvHsJS3
Epc3ltXl24nAYn7GrJJxC4qXpvKDKhVKMHnD1AFfrUC/hP6jqecJa11gqrca55JW
ff1OaBzVvWRR/y0y4w6Oi7aGqd3uvtgB1ogViTrcI3vzWhcnAy/cjct5u3faMInM
11HEQMB8kvAYBMgSlRqPgM0MbTIq51KQCwLK7rmG/4vMdUy4hVpPt/VEGDOYs9Lg
oHaw3Xlp/WbzZn4jdeilaulr5IEWDHzX+QlQTxF2vvBnEvHuhFQvrQiE70uLkUkl
eunBrlsf5QVFWaEdun74VI4hJYRcsj2/PHEJFZXz0zyIULDmwrkErXOD6t2qUkZD
3+nlFo112ZDMjj0GXKbTCxlKCA/4iBqUYRktXSjRq/7H6Cm5MAn0xxbeJkgqLm/L
yQJGiLVI38TiWx7bEnkA24ovgY/tl+mwhuRWw6G5xOr2tgPUInF7Xj2FkuWiln5m
avGywXdHeq3kL4g8HAMjTwTrBxEPc+dX+Be9SzIKMy1GYXkWunHtIAom1oCvog7y
ab6gK3M4C2x3EKNfXPxAyqwhvdPdWEclMKxBXHJt5sDd4ZTG5ICTXdTR4aPcEjxp
dThe8Tu4rQIfJ3KVqBQf0eDinsHWDqY6IwLRrlXe6Pajz9JbHAaFoAnA+j5m4IpP
8lPM8NHHEkMx/u5bzqxz5N2mqCIlE3XdhHf7CI+jDBGAhELaorKvfg1MdVvyqdtF
FdiFg4hqb0XxAOgbSbg17uhVPfohLoV//QIgLe9s9zSUKMkenmJAmICT8criIVWB
oXdMQeWu33eu93Zv4wrMyQQEM/hUsW1lKfUbK6gfjxA//QUCE2ymYmj/1VwFF6Wk
jViVc7h4oJeY1aKVeuj46criHK9t2t+TbJeQeuxeCxKA0ff50xhPkI0sOvoAR1ut
OHSDwOkc9ml2vNmgA3ijsBHD2C+5KTVxVnVTlrtngGUQzO4wPRiR8JaDbtK7VHiJ
XfeXPcaC3ZKvKB1VzqUMyzi5rn0l03eHYEMfrohuF/7lS5BTe/OtDIXLvoDbEsT0
wgQCKf3h5rf8O2ZVvbn/VBRoIwTAP72+UK1SSRQENuig/Zv6sf88j480A0O/xsHW
cJnFl/zqlRjMU8fYTFPgM9cpCNvnsL9lWIEU/UM3fxOTs4bX9Nq6Y1lJLv+6OGKd
juWQYkdhcB+a87ScCwTkRQpqGYhpPqYoPQOpcijtQPG66JILqvpr0Z6k6brOKbpi
K11CcCxyIzWQFMg+M/ZeATXk9LiVJgfoy0KQhROYHuL4Kl9stWEt6+wB7yMlRRgv
TxWHOjhsbsSHbzc6LFwJj9Iuvw0Hsp3c0UBLKVLBLPo+APLm7p41bKvjUhSc8H0s
R50cDUMwOtFiGSnRqRshROpBmWqFxn9OpYCiS6EVZiTEgSoWEiI43Xp3BXCHjuW0
eWDHw2nwmHEheGu86yaQV0M0mXW5bA81tI+oFLY4uwb5jb6dozi6bLCnAFtqwfgd
RSjFJRgbUjaroqEae2V59AswcuZApSN+JG5bG+PA4MOq1LF09LHHr3byzajzAKxn
WPzW4vu3w0AvixcPqhiEg9JcoG+uWLehAbJaEpy4nQoArKkVkb1ANC7EPxWQLMzN
5PMLjEaHrUjO2whlDgvTGPLCXKGe4T7uxFsK5+nOhuaV3KofFR/sZsnlmje7/e5r
AJ0fFmy8AthI2PNxhqzpHYJa0e4/SykZTODmkzwh/kRe6q2PFjpZVvBKRg9NyKI7
zPUXlkzbJqIgtlHTCEIRmz5WUcCeMCaQCj75dCRq/QPBNkz914WAgpeGXNBK5QUA
sOKOtwEyqAhoUDyd5rKqwDHI5X6ehM30pP6YN62l6JxJo8E5DhI5vF876R3KQ/K9
2VdWAwcwNBIGMhgjsgVRjLKgE/4QqHQGBoTVEF6T7Y50Ne+NIlcJWQb8vg4ZPWx6
OjcR4ICViGwvgE/PSalVU+k8jwDXEOqL+RH5veL2cnl3el4zFIA9nfaeTOanGGvN
ngC3W+TjXcqiUxronjrykJdMX0W+rfXtO+GpNcpclpJ+JOjR+r5m4OHOPQYvvHz5
iBnG6quPdOXvU7kf3a4WMcuyb3LMhoto+U20DiAOBDPNxQp0Ic7Dt9KSdNMws9ah
KUxcONdSzRZJgjPZvi6H930t2Ik58mVshTwMtYXanWlAl3g8zP3FbaRi+tbmdDdH
e83qiVjrvMlcFH1KcytWX3B10y4LFI6lLlcm/iPMfO7uJLkSg/TAso6iOgkmAB8O
TrGWCM5ldVkac/jHFtMZvypWm0QyenRi6lQiUw9v3Nn/PgdVwINmbJsj+1cH0ziE
d22CpviUZQ0x85Vr5Zzscn9jZZJfqKbRqvV8cQuMBYOCB2GE4n3tohgi52lqMXZb
yrKGHjCMNqS+Bngo7Wmyjs/D/rYuBKyCG7aRQJ0MT/NZROnkcGz8mC9gEHqDOttK
k30pBCaDrOEUktEdUzQjOP5QCYsGEaLD+9y4ITg+5z5KBGn9qexgWIIThMSdwHcP
Uhujg9NbdXj4xRcAhmR1bFC9jJ4gCEhSLijGpIpl82lewoDTjx9TvrYEKZGeVess
CXUfkrgV/YuBzXCe6y8D80sAG+9OBGcuBVQpKr1nF5t/vmJgEXtJNuEHA9DVC5fB
kObOcOFloOyFYFm1xmn0c6h2xvJAkfY0lyh6K3D7hzFwFyNewa0byxg31ikubkxN
CjX3Vx4eyA8aVA8SPiQuXcrHZUAqb+RCOirKqQr1VnwiKoKAADDD24BstN4VpISR
uE+hvOG+JFmJNlv/4hvAXzzDtM+bzcpoQyNx57KDnhmxg/Ko17DtGG/ypoIzhfDZ
dxuxZgILrHL6SEMWk3JYeWrF3WURloQtlGU46rRzww4y6/YZfM7IV/YqQOJkg96n
UcZaDhflsO321eDJjh/ammghJUNYSUWu5wQxOC05Eb7SsmREFkM6gjP2Vj2nwXp7
FdbLIGxxEIyYLfAoOj2gnckbhlJQ1Jpysf+pZoY1zq3LStApghrFjEK9UiuZgqAm
T6ccAEUoWF5F0XPIb7bQ9/ZUAF80Iqb7A1/NYjvVrkQkW6A33NJx6lG8RXEXrxiu
+/xXDvuwfbmXRsJt968AqxdJU2jUIW0FC59Zx3z+zs8m9fi7uTSybFvaTRwr+YMz
MfGjUXuyvL59zJIgUtINbNQ4pd6ZWVVZEzfDQZjjJmNEN9iyv1yvk9+Zz8M3lnIL
m8wbHTihc8tONb17XFnYCnUJ8w+Ijv99Kh8e52MViPTPmgSErLIIZkDyAcwqeK0f
IohnepuZXvUKGLA+omy8udppiYeiMaPCniFfqa0mID3c6Hu7q0h4TDBbYUVtl5ci
ZM89SVDNvSOJ1YEPVxSPNaj2+P3u8F/eclt3EI1vmxxIlKVtLE4SNCYm3wEtLrjX
SGwMqeNkrZOoF7/3sP5Qpu1E+3eMiC7DtO/Klyfe5HNumsn+PXM0ODLzMMGIW+ES
D1K44Xk5ivlxMWSL7Xmf2gBPJX+9QO38SIE13+01Qwv8iA+CCBz8q5BFtZs2VH6F
gIcVDkQLJ3BB96PXnxXrPx7QI7Ckwn+mwUqmdcuopiUnikbie/DAJWe4uVzFGN5P
oYDk8fkz6OZhyQVK6ejQCAEBDlllY1I2HjIEQf+aaCck3uQ1OTcNHjLPYC5GhJv/
4LxHHGnFKlufiq0nDo6i2RJO686CITzXVMLyiVMKfdStpbzKWrzZRQsu0t1AWI+g
IcEWUeA5ARH6qPTRL8vWkw6spkkOSVqYPn07AKLLFK3qrqgP8tq183cxs3d9G1oI
uIqqxq/TNQWw8WGL26Tdz7lSolcHNaoKgQo+FqaLZ9WdZRFGdORwgIA+DEFGZf2D
8b3pBT4se6ShWQT4oe8ZR/3pEAkyvV2dKEYgtFPS6Vxj0MMSBFunlzdTB+S36GoP
uu+bGLFQZllD7a8y87VJj5Rn4J15h53ksHOhB7GDHL/noxJ/nMp947ZyWyRz2EMK
v5TtqLVLhOq9Vrl8oCanrN2Ljq6UXa19/5nkLOapTjsBEuFgU7+XdMvdgyCq1ieg
DoEg5LmPLvbZoT2spmdYn5sSmcTki/8xaB5wlOLPbdW4R3hk0kmJPuh44fFC88g9
O1Ck86d8fsb5M+X37ohHZ43DmRPIGOByI1cwhcqN0/kBWaWgLFdzhqKjaY+8dqHn
BAdxKCrd7WU2Cq9QQqSXCgzZQtLTSlcKIhi6ZUfn7YYnQMkTNQNBJkUmshc38KK5
eYZNdQc9Vg0+jv8S5WXyAuLUjJFeUVubtpRNINWUZ+PqMrwJEdLpcLuFxgSALmtu
+1wfGYOcRNDAu8raGLYWFGXVsHIgCGT5VhT6YjTlJyRK3Gq3xdpJdknvLPckcjeB
FNxxqXtYSvCa8621IHrB+Glhrt4tvoCJqduuAfrE0IQGvfIzzMfvpYEcc5j8DrMw
TVKgkYAUNyklVeU3MxUPj7r8I3sffwGgEjxSF+xUyiUPn2hU+uf4ixKyTMX470qG
iB1hIO8eSK47mnJImBO1rnTGyRTt/OUmrz1f49PfI8pnYWodaIovU12y8tPGRp5w
Aif1MF7JQh9Wqdlmvgm1U1eDKf4tacC31un3WUmzYMnrMJDry4vMvjLs/KybGxC1
hqJHXlPJzoFpeJ3mtVnRqXcWuTFrXW/fci/8MGW+B1qTYMbIRB4/k9q1lR5mbugL
xMGa/92zUG7S56mcC0nx+o4CAH9wTPMoLcG3TiOOMRR/DzkTOGs1kIFe/YYlEWh5
ED29vbxrOMZh2tKtiACkw4NVxJhOOpJpk0EI5db4Fgk0W9PVfe9gMIhJ7IDWU1iD
JLAOnXEkpjadRyOTLFH4pdSYJhMMER6YRJ5MwWF6X2gJyre0jE7yeo+8p/ARUcs3
3pVnYPba5jeqCT79sTvAZ5GluFvcDg+Z40xgU9nDcQp1kdsMxlhvxJq7SjiZOf0v
w6L0H2XojUgzIYsqs1b99Zaepv7SLiSuFxIUFP9GYfCzHDqr73zt53R+iz1sNz6I
9bDV1lH9hceszQGdmJNySwK/vhgVWP3oG261Bv4l34VDcszZ89lmoYc/BQ9Dki+n
qGB5KhVEVuXEEBobxGHxwO+t8w5H8l9r2WsSQlwk6j4OOJoQ6TwRDjQRON81BNOF
rHpgEpQKtvaMMXrq/Ryl6W+A2Eme/0EE37LA30DyRUceGpwqa9wPdShMTmQSS7vx
vD1LArnHua1iys7KewnItSmnDMm2cRX5esg1qDynJpUKtfh7y7f+BaVrhT4fphir
ue9vVd/atGmAy/XLIa1UzbrPK4jV+E4zcle8EOdmwanZ69IvYpZmy4hoG2+AbuLb
nhDEN6F0vsfOteeo/Bi+l1i8FQSS6JW+/IioldQzYPEpLDKVri8f+ghgr09EAcAc
204D6GucUcBFQtQ4r8VpdgCDjYqCSwcYmMXBP0YCi66M6JTM9r1vF7MaKEuvP9ZX
nX+Rbx7MTjrc6SBvps12BOjJdxM4ICcrwxQYFYb+lVN8xZwddCxkHbX1efnFjZj5
rG8VuLENun9qA5t69nQbOWYka3Nx7LseA8VNr9Qncs50zp5mhI8X6Th5t50fbkI/
okg4QDXkGAk8TIez1g2R1MmBjXqKSOXPLsw6RVw2GWL//f/dWcYhLhnJndPcpwwF
efxb87+NC+TCNqE05Sjm8kc6oxqjkOCihMEGuVJ/ft/XWrluKNx9LvKJ6KU7gsi7
/wVG73+uihAhtMCgNrv6QxALu5Mlx7TVdvtrm5k7sH6iYuVQhi7Pz0fETExu6JKp
7emUKU+3ZvlXU1IT+sCDUbk55CQpU0iKz2HbE3Q8Fy1JaXntjKDGuVFP0ekYevv2
iFWHOySubHJirWlFN6sIwsibISX92nZwCF5/ZFIqUonasblZDUfGgVPAmWLrdpOi
YVwYShvGvBzD2OoX5D1ECDidQ8PZOm4VSgpSAwmSDVb7E4EaQc5QsE6/oHJX4VMU
Nk9Bv6uQiwEOmdt+UQlre2gv3/1l/qksA5pKGr/bxhJMm0Eg3gl9xO/ZzvlkRIWQ
sVT8j3c1qPReDDN/T1jOpJZR5ChO1U1Oro31kJ8wThmYgyESrdUUc3XDi5AIGn8R
xEcgXxUoHDBSpr0I2y3NzABppK9pNMPUbRdfwP8X8XQGhc19Fe8HgqgMOW5yp0nE
emnIMfcLDJdHSbfXw8pQtAXEmDpdrVvuIe+oscw357Wn3Zkx07P2nnr/AgHZnhBP
IDgRjz/NGK3cMSPDqOhJsji3xLaXm0jx441B/OIETQ7ZviChmHKWduTY5z2qPvqR
EN02lrW24tbA3EQYV46A6BbgvNMiyHjuLRXMgix4soHFXFIe2iMneEc7Bl3OhiPa
OqQRnkpQJ22u1QVW5ARz+CAIrkf5R7q4hIcVbavte7vLfOiE8rKT5u2UXOdF8cPd
ebxMXu6Lbe6RpjznzM0T2lkHtLo3RusPAT4LSRyH43BUlv4PQOYqDocyUWksF6Pg
udMtQg3i2koGFRm9Tq0hp8jouOHb5t6NnpD9ayMpWpsq3dTw81Ok3S+fgoEwJ+OR
qrh4R7bO6R64xdiuWI6IenuwBiKCFIF5vaYSFeETZSk3a27B4hMiormMpykexz8v
2YSu1rU5xbwoYfS10q0t8qg7gxyMpzsq2h5Vv6wfrUVx+EAA9LTeR/QqyfhUCmRT
PyjSs06awywgq2tmmarT1j2vnzX60T8QbS21E/NMbLls1AgwUtyM6eL5LvL66miS
VpTqr4cGUSp/op/Z5UgCRAiZ27Z+JespSuOh8mKMbpKZBNloj3dqZMGS5q3rMgC5
WY0D8rbUv+pelO0ex3hwMLfSX2vTiy0sZj6R1DNh9ned/en41xyQp010VmZbyeoU
crZa6Nqg2hN/YzcTbU/uz5uev/u77MdRfvEREJ4G7yPUvH/GerI/5lR5CvOpTSg+
tEWFMo8kUJlR9DbB2Z2vHCvTP5p1M5L0YfplBSpjZoTNASyuNquT0TWt2p9Jg+v0
NeQVyLqKFOJ5+Un8NUDAKjPXzkQU1jqK3vHTeGSD7eemaN+mvMdhHOQlgceuoTKq
wFBXZSSSyZSlCz4xfDIP+yPK8BQ7AVvGbEDvgdK1KmAm/Or1NWZCcm6NTzpp1pFk
sdGRzl1Lth+QtBGbDUXZfNWn/Q/WFDdDVZQMrzXacVurTWHe5EARZ/amV8My3tbI
zmAGTrUMWMDVStV2zVn+mlD6D9X/0/+jlbtmhpRigNpUz49gWzVdVNGaLSnwvzDk
3UZt5tlnqO40JcwuvJVPAQRTgVQMkcOk20+wAahteFWalNheFXe5SmrIVV4muko9
frptVQ0Ib2T9VAqhKHRna5Q3PUJW8paPkwSTPzqGumHzpzLjGFYatLgCOwi4bv3T
Fyl9iFs5YE8JTDh+F7BQyEObN4iwYLagyMt0YSKicpGf9frW8hYm8YSFUelvu5Wr
H0d6Nhzp2KsosP0VeVWb+3jRd3JYHJkgpB/MdJ/kFct/oeeyVw+pwqzVvZgXYur3
bdMp1Wh+MNJFeo+9+dNJfP7FBHQ4wjro0Opj13pwtkmkvCCM7qgN/vI5PsuhXLSb
t7vWqpIMmmedYetXauhX9vYArSXaR9zNVWa9Np2ozcCGdHR2vAU8aYILfmJLb3TC
Fb+EhWZTeyKiBx3zuIVdmQKjZ3J4g1M+lUuIQ+Vk2y6W6INKtwydKTlOHKpZM2Xs
gFuSRrui0q1CWJnLhz54zRjTZ1ho8FvvKbaR6B+mDKDrU+pcwc4NUmjiaYKZKbT2
Mri8zqHbbB4la25WnKX9XB5s9b9h5bfbKxVz6iaF38OylV2fXwM6F5Rtf767YOfw
sVmNI8muzZhohN8jED3As4V3cU/STUMqApeTafuIiUcJNOf38wJJuETGVWPLQvDM
lLRGOB6gH7UoWYLeOWex2PfjGsX869n8SBZlVGwGUqnBdEnyYACCw2xMn95rx96P
WZu+1gUmqpYSST+tIRTyHs7YT7B0DgCuZDcvkmPphjGDnvlVDzaAyELEh5tnR3k0
KU3EotFMOskZX+MmVZjQOYAvev8fJ1yVVlImn5hx3amWbmBRuc5vlLj34ieODX+I
SS1P4kCQthCJD9l89eTBfNK3OGw3Vb9Di/2Wtv5sA9sFWTBAFbKs36TKZGU/1zh+
eWCNLaIHtu2+butjcfNAGrS9qB8lzeZFlNiDIMFs0K8V6QgsvG/sAzKf9kanXxTC
TtmTRyFW7izLGtyvCOxsUZS2dpludo7/AA6K9LJu5rg3BWoctJZCjthVu/fFUbF/
b52QWyfpJuJVAvibRXSw3xk5O3oLgbo4IYxV13ZVaZugRb907uLLnS4W9X4YUOMT
zA5rR1Rjf6++RwgHdJrNKT2WhTAJ/Nm+zBJgz0kqaFVZkYAoeHcGmwp3ch/6P5un
5sUZeo9fk241vwv+wwVA81o2y58Jcs0/w5k5Xv7NmEMzBw26XrkEOP/AvigyDocr
Rp6hBbuGjAESUTUCQBg5yTVI4vdttpuE2uaquNNeLzfEV7h9fJ6uiMxhYyr9q4jF
OCwWTb+BajjY6cSodaLhUvE7hh3giLUOsEhUJdLTrYKeNflSz8EhyhsZNdvNk42m
n80gaG0urdFZ0e02bbM0v9tB4XaQ5v2NPz90Zr03hUUogo697ccuI9/8e9Bd4Z7W
e4hhFxKTaPQIZlts0QIBJpl4LD9M5MwrK6E6Vwrn/uQhmcaNzuHGYfJnCZ7a3YX5
Qm8Zwr/LzaGLX8HDAdbbiY9UeyfilRFAth4QvZ0W5lQe9OcZDlyx5cFaya6jc5XD
XFY0ib7OBuRyvtJZJkwlJVnwTAwjuss+/594T7QwbnAUAQCJmdAcMDtwbIzPjCMw
xJ1yiXT/yB+BvJ31ZiX9jQDDJmfll1wOfQjE8ZpmaFzQL+cQYZDR8B8B+yLiHlJg
51QzuKWGaSeZHl9vYfRalNFpIqT4dz9f6yTLZHThgskZn+6/1B9QVDVL7aCSfWHH
o5mo35EB9+Xv8rXoX+/QGhmiYFD9IOgAfVVEIlkfDl4Nnu6lRDiBiz1GITXrd29c
zDHPvzP8Nj6xyx1+QJzeU5X/FnHVqALXY7RLGi6ldPxDwqXq1+wGZWGC1Ghpl15y
uQCMwIcu6tCSllW8dCck/D8PSNVx0Gzq03yZCV9ivhoCjUUE85e9flkjEM15F5tw
wpZbUPPke1E0CoOWGfiqUmqsUFytvEa3OBKLu+bGPdUZB7pGwIsDXDN2DDJOgxpo
tiJmhqviWkKVX9M4Ea3+7WBHaiQ47Ho2hmhYySDZEQBhq4XnCzFhNsocPXaEMpkv
qb8X0wa7jGw64o0/R3UvuLXowv9VHoC5t5HveOP2oRWzhxOtjBK6tzWLCva5oXlL
YfMIME/WwgXOwPj7rsbakNMLdHjD/GfysRMhkM+3hgz/TTfOWT7By3XQHRL+Rt8t
aqcEEvXFAxzaQ8+74WGTbxviskoyL/6JUSgK3wcj8lYldo2qOOkVq9SB/oqvEQgm
sSsff/SiVFULbYVhI1mbOKbx5TYW7R6cUQMUSvJ5kiczT2RPxwYNT00zIpByD97t
NFBWLvwQQ1lW4CnscZJbQzRUKc01V2e47PD5R0jI9rEL2247oh1EUBBUfoXn9t//
b7mKmlwuI0dcwAkN017JhtSn/xmkxLxSiuY+ma1ndgkOLGeUruhThtLtDp44bYBk
/SLADL7Z2EEz+OtTcj+lHV6SQuQUoJ+cj+aab9HdPqxYXH4TN+erbRI/L6ASVrN7
saYatYHe6wn5XwaeQLMtjVoOl+PwKUMS/7xNjN7dcAS3oVX8D9M4Qa+gJMxV11RZ
gyIRY2zVtCT8MukNYH+H6wxiGATaGFGUlkyvq3EB5WteZbskJnNRXErrzT4gRZSD
GXScGyZP4zboMrp8poKrx89ES9MxYDxp6OtEDSyxGUwcedsEZJalmYYCW1tN3UUs
pWTCK2KPwWG2s2TtYNa+g9XJr2kxc65hlEFxjXjNUGN66SgDq/C0lF4QC2A8T5H3
rvyhKBkgvhLOov6vkMlMDR4f/dUMLxOhsWL295IkaPuW73CbaF+MfJkNXTKMbJs2
y0BcLIlwdatsUdFzoIh4xt45FbFjZX6ddGhR+wWT4CrIMKdLXWiuqvhCpLkBEReU
35rD8yQTZQn5aH7eB/xDv2CBmcw/6TVwnBgKfPZmV7OK1r56F+3Fq1HFxXiv9MxZ
B7UjL6pWDAFOhx6GneqV8j0mh4EAyAK82khAGxJLurvG4LEZ8ooVIbPquwFKgekS
UF3xpIMbqEdUE3g79uFYNjxZSXx+UwaSoExcTeA6jH0AvZdLQ9Y94xaEDSTmtKYB
GwxiZAfbPSUWnOTDrMiiszTvgVHQz2eoQ82acGOwLXZ8/ruaPp57iZrb/k2qWqej
pw3C753Q+TPyQRUSKRl2YtKrgS/dyHQ8u5lln9BgTu+6pSNSKnSWw/+biEdT5iaz
LkDuSWJpIpndknc5fL+Cj1eWB54L9MAhYysAV5obC8grYMeKCrgUNNRbmIcNQDl+
kxuKAC6UQAkS2+01wKuBU/F3EQla38h4AOf6AHF/lpap4uCFii/03NYRY+JikGtT
scXVrS4U8TlCzGMGNXCgM0/cQmPGwcQgq1kKFpH7bqgMTwlGzxcceNOmE7yEMFAp
dEkoBsXx7QnQOTD54+4a22gAoyE040R0NKEi5HfHxua2XpuSuCiIq+u2IqJpdjq2
lxtu2aSXXVJRw7uHpq/l660/UYDCCQgHEgD/u0S2V9yUHoeUz39kayqoy33tQq6j
xDI6zpDDpAaCgCrAKonVyYiN29VbidUCh2ouqs5f51kmIbn0BBNCoN0Xikq6gGjE
Z9nmodMbd2aoP4b4NJyKm3pW2RNb1hroArYJ/AiOeGDarQCe/pBl0wR4Yq0QDwrU
+AHQq6Iieq8YV03zuUIByoRYZ5z9dXRoW1fdYmycNrIoj9V0r5RqBvdl6gM5Gnbb
VeBkq3HO0rEARw0HBMiqDH1xVQ7+xIakobbDNUJ7YhVICUodzCD0/2sT+BCNC+mi
EdljDspEX4X8UXZ9oMv73gsDuUPJX/UxS5mM+nKJjewIMS1eHJLvWY5E3MQikK9x
3uQWqEPHoVkfKJuI7XuD7aex4Ckhq7+rjIVunNG987UX/W8e+Kq8YZ8BOX0sBTgM
5CzMLNU3yEi+Wf+eu1hx212wPS1jOk+++DrZbkj+5+9pN5FFs9m47lRbRuKvb/2b
O5NCSURjcBOuvZc5u72NhnKv8vPM6yN9Pg+QivDIF6DQ4jTOHenfUvbJYLaLtQzG
OyVXV6cn9eywAPD8rSU6WsA99S2T24sEwcBjxQE6WSh7ITYASNa97RPMDW9+PbHO
AKvJbh34vhxSTFveoI9OrrvhnGEaDZQgJqxArpR7Negw7eBxZ03Uey5NG/tvnlSh
3wk/Z/pCwf2Ufmj6iKoZvZTaVf1lWSUjxcRhwnJ95+9Xni8iIbyZbVdveYFk0OTN
G46tdUKklHzyaVJ/1shAKP1scj40obGckkOz1qiYboBUEsCknR4TixwtfpLS2Bet
cZRU0OGVRjxvmcbmstvpZFADJVz3rDEYBBtVUPPMZJFGGsBogp5ZK1bA/CovV8Dq
YmdASOzI++8/wSePvJpl/ANzd7+KKG8J8IoJSNRyvbKsN8ifJIekeQfEcDO97tdg
7AEFzFvJ9u5M1DDOWqawWwEae3bmBX1/YIbF7CyWrohy21VxxgneDI3ohWDKzEWf
y5GC+tcsI1OvTig/ZHKebTEyGYqvj27v2jdM/YXdyAk8rZhQ/VBTWTT9zvknvBic
L9h8LmUQhIXMUljUffq9a0zy0KwaGuw7TI64vv9yQwE/WABS6scvwcoAwRuM1vmb
EhgzfFU8zhkFYIMY84QJf/0hyguzW59AJPQKShPlydyTOlI/OqTLTRGU1Drdg7vV
LS9y1nJkzbGYUJfUd/t9VliLFUEnXMcvCdRmcdkMNK4KM5Fjptqt8/49D1+WQiSk
rJqNpF3mcHXEATQHziMgyRwf5lRCiOeum3UPe825t+jb0rI8/RJHnwOxniqDG9x3
/pohI53vjQh2nQBP+dnQwKBS7BFOB4mBSfn1ASRCU5/Mttl61t7NOGRkV//zoWg3
aHJ6JdccCFC0Kct+6UyHJgiCIVUATTeSlhF9aE+IVbL9y7ApfZ/78HZ+g/I3hxxp
OM6P4HteElciCoEYoW3+or46nSm19ZL7CzNdZz+SrwUgujIPsAKnoQGB6RmkU8p8
xzr7MzUvWFU2w4LUwplde/VOAxC1heE5urpN/q//p3xTRXc/Z6XvoY86z49PtrML
siLE0JXsVgDbD5ZClVShUl48YX4RF9EZ3Q9eNXcuCkv+/q9wQutXa1318GT70BmP
VcRgJ3FZuymhDglSg63HJSVIYKYPQqDvY36xnQxMF0nOxSifjvzBmmSgIFHa9jIZ
Rseg2g9YvNP17QFkg2bVzZYCZMFC1PMw+sf/J1gIP9tmaIjBni3PZbKTLkOb+fAw
d9vFe1mx/T1E9q+VCeRGQBLcpsntm/dQYZVFFtZrxQephq0lMX4zfvG93/kHGySl
SGNNIVIOy2eGtPxp40Wcm46kDLKmBhZFVpnai7kj6BDLU6nqgSv0wYt1acvX7T+Y
FPRdWxnxA8gzsNpf66rc2mZAjuYVmaRBSqhNwYXCyxk18vrYp+dQ8AC9Cez0STR/
pOejwVCi9K1y3xp9WpvXCX5NvZaLCNRLtqn8djldv5/54lOIUXSzZGhRAm8u8Sc5
DUsF960rt6Xq1LU8RR7A9GU7ifRnKFD2wuqT8z10L8/JiVvnlyNUXLich7H1BOkP
iIaOQLq/Sb4GVWMlIEyv4jcyoRQ9TXyAluDMwNBspYUqTLZETEow4TFJu8QMynzw
LBhfXw1BC3D1qAKz8m1hC2usX//a+l3/LDNjQyUf0bYRFLV23OgQRFqq37iYs4RS
TQgMVvBUUd3aV+2ZzvD0EFLn4dSI/nLb7k4QJCozL4JcCgvCVVfIQSDAEIWzXYjj
fe/9qVbWaLeYZK3HK45motFEWrevPQ4ZEm8qNzHQ6GPMI9sG/y8p6iRhMCcbAwC6
yhd6Ul00QDJNKjbke4r0NRfUP72NhstZCKKXBySsw8RlFthZxk6S/IQH37gFtXZu
5u9LrQxz1I5XcJ6F+yWse/n7eGUQObj/043A50K3Of7CpYvFfsNS2Hg60Jwx1N8m
aTeE8J1BW8hmJb2koXc52W52wU0oTeSq5BIiVjZYwXcGyc2HOnVLUspl5rwE/Vmk
DW6rKKMBxprd4y9rIzZpcXGirxCxEPYSWrl51LJzH8PlRVBSIQsQzqgqyh+ne3wP
DDQWIapgj3+cVcT+zMjXLKNYrq8I4rRCUetuetYdpV76tRxnpH5yZC8/FQeGKNsC
+xf1cKBw8ZCVm3qAWNpGxBdPmF6g8GvEAGldntUfbQpHaP339n1OHU5PiqnJbdYS
cEaIoYwKoLPk0ePpfJ4WAMQbqVuiMa5Bl4jL3cygcE+IZixosoyE5UgF0N8M2tAq
DturnDjK/W7imKU1ndl4g4BDvwaehA9Zx7DkNap5Q7wvzIazQGQlU6lJCtRd/76j
LFd8V3KxTmHoxs0SZjt/NdkeT2OXuoZToionYg4VS307uXTBTJN6KJB59Qvi5SpL
adaQd6MXz+aGaNE9rdPiBUanLxpy5mjW7q2YtZdpQxKoipYUh+Rm/4W5EApofl5i
P059cS0DoC2TmBBs+TBwVmchE9D7TWpDgjsZh0kAtqlgv4+lTRWEYEt48314mI2R
ua3q7vh9s71JqgJFcUwSUFQB3sktJ/tcAjk7Zm5ArsrggkcBSJhvQRbtt0yjlUQ2
dsmvFY8YGeJqxZqddulUCufIyrpf+HFkSS38F33109MhK41njQjpQRU+xd3Y9w+g
dTVxpDPdkPn1VuyEXnvqQPmLdM4EDVNYwS110KtX0PHi/ys8rxqJlDjvaUnf6Ns0
BRFu5QYeG8b1bl7U6xfGvNvYv+2H4K13N9kAOMkeVewqlk5Id2jB/k9L8fBOfos9
84FZxCaOX5ixhDNuDtlaavhINJCz7/xladUseF+9DDBYM9wBALplJ6dlHwSftgTW
iwGWl17DR7n5UmNUzScKSwyJmGRKdM1UWJoB+1TAd0wEHlm5+A8XYgS4F1vRQgQt
cc90vVY8hJMI8SNsRGsMlCrImRWFtlAwAkIAsHTxIacn7uPykRNkqcDEPCHJLqTj
syqhGtqvOC+NZyUv4DmS4IfbTtLISm7oMkvVlo60dr7yZ/d+HFc7HuA8V6tNEQHx
CuVOzPmBzsB7lXpMj/xsLCUe0huB0JIQBO12D/jiYHzT4gM7cYQglfN6+FwFDy6Y
h4c1MjigQsxewhty/PKHAoxPBK3k9qNWr/KU85GEIx2bEOxl/3o7iRSn7OH/gQz+
Y1b5vDe+hdW3dME/E/J5nxwWFbCnT3/Ne4d0qiFnsGjAGWpDtTvZfb8wx8MlbNpd
iRtqMcpTSQO90iUbw0TzQuas3tnhMG9RpJUWgS8D88Z+Docsm6oBTswVmdRrtu0h
FFBAn9k4FAkWpYd0+peGqgyEGKq14D7C2txiFs6g36YeyMaMq9IEhTIxGGzB63k8
zvL0uFQalogyDT55w7TbPBckMYVkUdlH1xDTPUiK8teIoq5azA8JxE5EvJX9PMEy
SmOuTZaG/3CkeBiigithi+jRXpB+SJTeevPSua5ChgCLdZhRUCdME7Wg/clNc/hr
WOW2Aa/7nhSGpPLeGLDzMQYxOkK7dCYHHtDkkyuvbb5Y2HmM4pT33TJk9UZ+0ntd
XlCVfmqoxIUads52ApB2vjz8si+u4QyKRsLzNaYiXwVEJU9gmXFAIknrHgnRhnO1
WNpQnDUVSz2HNEFWzDJcOT036y6G9dFH0g3stdvenrC/M/RWzuMHa3y8Zi9foNFW
/2Pq9mjAychjGCbAQ1Dikzj4LG1RIzk+EpbomJAUwxXwTzenYl+/15xZmWiN4MuL
ItlDTQGCP4UfJo5wMM2nTpm9mOq6Mg8ooN7AxNJvMuEicaVJMnwCo1q1Np3EmPOd
7vsOvddxDSPcZsmRS7Yw7ZX5dFg20UHgkiFazdYFRBB77at8j5TwhH6tIW8tq9Ic
M5rWM9gXJM14+48A11vrKCjm+rMSEpt8JpdO5CChmc3gb7W+UusjriWJ9H1dCJ1a
frsl5lfhh/vRVkSfxC7EyLo97w0rFopK8VcTgCmDp0kCPatgyufZomjxaTA1uDuG
eJPveB4ixEkWwxmtwnYzJvUVHckmT02gbcIfGoGCc6hpQ8qArQohHGQTTr9zMTwY
0UNIDHfIv3bAhl6Wbs0eBjEhB52EMUNy60OduylrKmwrRw4s11ZmJNAFWEDuyY0O
LOaRplICK+NMHy7EuRA/j1T+3nwKlhoU7JAbkyXPoX5kpd6iLChmV7dNVsJNCPOU
cpVeVSW4b3EPZuW0t3xOeqep++OUkiMyQ6LiRUPq/g4jV61xweE0NJcZu3kEQHft
sv6YwJEvxYzrAVLDips6SVsJ1aA2AwX0jMyyO3iwu7ulmE5xeceFBlt1eruLm4C7
/eD3datiQHRJBp2c1K2+hESyT3TFu1yIvQvegjQLr09cLd9CSVzpDmT9Au6KOkHX
wLRGRu6cMhdGULI5ehAy9v7Ik0uW+9Ua2kmb+vS0zGyG0DbF87sKAM1gnu6aWSbr
0S2PZ4DQn/hiO2c6thLZ6L6BISmUugx3sYase7b9rEWKsbH6tMPeg2egFBZcO57q
1n87wjMtOO45Ev0sTcPHAalO51snNkki/sIpH5dCdpeQoRrsad1lVKTe4AidvDHh
N6q0Tr2Nz7+1tfCppxoXEnAND2AKc0+C921LbAu/C8jU0PeZmYnNoHAmjicDhLWl
RVyUq7pVPjqnc1ZVfhHrlTphnH6q1arq5h34dbwU4sAzn4A4HxozCGvY08QSWMtQ
m2V0y/ztjLO33AfG9Ew+pix7BCbFMqAp5wimN6jwoWE0GCEJvHToFlYvbSIxlzQ0
37ODjZfOcduqeOCQE24J5yz5WVQTOkZq5t7qiWWjK1WVj+nFyZUFGejhaxC+7zTe
/n1rzYsrgrMS5/T7dMM/DZtJEWjXkdCzf+ipFKZ3uzRyeFTw9cF0RATk98PFTvZ5
qNOt80GCaBcLdgPEXflW+sTrnqAXDxl4tEGvmw16kQfWaiF1f8v9whlDFwASIXXy
1wIBKLSHinUvKZO3Iwni9968zP5u0hRvjOp1ccydpr4GkDMpUjKhrjIwkx2wjF2X
aU898G8RtpAabqf08AU6wIJOl9WpJcGJ4hUkcqAoM1yf6UlM7EnQsfAbN00S2F/w
nSoEtyoORQgpf/CXBMgg7Y3lU9iShRTIPTHckBd+6bH/RzNxr0Adyc7nmudIC7x1
p1iH8q6+6xLveIIgLO7RbM87NbvPDgHgO04PRdBQ9d44PbdJwjwuzFFe5lxXTM34
I8NnSST24eE31WCJXXnPBjj5Y4kqIEUw2GtbmGvB/GfdiixBQpEgricDrp8wrY3n
MsAttq/dNnuH9PvIOreqPyrOC2ChQSMSe8MhMWG5m4fWfXYPTyE7F1cWQGHTR3rz
88NrtbRfJJ268C0MQHDlel5/N0vxGkfBzZ1rKoeHWjMwbcJcguzCMixJizuVsphk
uIsBYYV8G/Bdrh2vJemX3X5H9UO0akalHFGoF5/Ye4mPL83zaMfcG2xlrfEkOl/l
8QRjB8G2H+w7c7HCA7Dimdw5pbrURjLSX6HeJrOlTZ6U9FJcybiwQV4X8ssquVPS
0QxcyZezdaSpZ3fMkTd1bj4xdPEJ0m+YREiSVW8m+c9OK56AQwy0xMUT7KRIpx3C
gJY1mWx2X0zdAmAmKcO414ztCc3jZqj9LjoOMT9hfqjy8vyh88Z6tYMHnGkxykDX
PdIA3ymY1TpbF0nF269RZBVvxWeDGnNBOMMWCF8OcZaqIAo13fb9r/A8cPZ3TU8C
s2TCetfvVVlA6OD2xAiEmVRjWjn4SqdiAriloxdnRRK++09TH92NXcap5ddB/mpM
0P1T2BbsmJpnb2aFX6W41l514EiSXcuB6N298uBqX3D10P+VASBzbuo/7/XL+Nw1
xsc+bGCjKTLzMSlWMMLIKkijGExHF6VlDB2xB0k5fajUJ3SjjMrjGtXMObRmAzxy
t5BdUfri0Vby4fr2KQMSPIIuTG67CtDlY0CW1bdj4O0g79I0C8uRn9svIQwZ2oIi
JolY8PVxiBTRu2QZ0AsCLG6m+5/sj6ksXhD8Sd3noVlrh7BCYi2u8ss0DcPQsEKZ
aLfsNgpkik3BVdDq0nwbYT8XJCb9f2GSRPx8tj/QFn6Vd07XfvVxBBVKIUruUOtY
Tc7NgTx5CQEXjfw2LyOir8xMAJNhB/38P94wkPgG6DZm3appGOZs6KcizsdOQ6DS
2Y1kkgIQpNoGVK5FXXCuz1tuljTJZOTMg3tTteb7gWxzNFhdu+u4t5q1nlcL5fDF
FUgtd99mNyTiGTvMM37u7zOeanRyPr3C+HnU/ESvHJIe42QrkkPz+w+WIO4/4MWZ
7F1u929hnKKFTKQuVEgxF4PZKrwYIOu2pTi3jahJEYmTdsN/DBZm2k0Ns+2QdTuK
p6YMJwOFCK2GuU/3Ic2T2pReRdivMyv497ZWrnr5b5SvfAxfO0I2aQy6geHzg2vy
XfUpRbs9M1Bth4fK3E9lLFZcCd2SJNZGwN5VDuXCu8kvfolHBG/AsAzqi8IJwMjW
KQla7nVcN00EZ5bfjVJQ0FP6tINtgwlDLSvSZ9jh/MO3KzfaJ9wo+ee2X5+Y++Jl
YrdH9o4p6lXXAs+c4Mpf9KSlMX0M16y72ii6yhKsN6pSu6p71Y7FLQWPGeAiHBb2
suw/IwnAPg3RwkyqLrNpgho44DEprxpLycdL395DOXjY7SA950WDpa3mGuJNXdUQ
DI3QOUpq38k9T365B9epl1v1BEjy2m1wNZNQLEoYof+uvKoGqJCAyWDRDkvfPXmI
vWqXEVWxr7PQG3g1YXD8YVaLjsFFY10nGLuwNnhGsN3WBAfJ1/cSGfAA9tHBaQ9C
Pa5kmlnFtMReYtP6i5eKAu0uehbJCpPIasKGOim0YVrj2x+AIEyxiq8mrYhJczNH
tHqPx46qOMKlowS0K+X4a7xXD63BV3NzrsHo2FMWtcHhkrjWpENWe1dSjThGTrZF
DQeujLKBdYjcBhqfn+O/5ZffUgOqIGs3OdZtNJAA/dBl5BAeF3FYCBTlT0M5P78u
mYl8Kb1GdzlnCh0RAvfGHAqt9cjJ4+K0sQTthP0gAgjTWrZLhK4Eqf8ksq1u6qzH
XgpZ52NNFoO8QdeqnL73WrBhL0MziSEc/Ox6IhUukTr1uae+/EUp0f+yzEiDHMRU
gIcdAFRtS+2Djd3F9Ae4zTabcx3AjtRvWNJCxftgRl/q6Qx5vlVK5yh3jlz2l20O
ZT9sQtvFlYDr/Q5/asnwH5blAQDAf6jthVmcI5Dm4hseRQmxScLRcXCeP9u1u8DH
e8S9ym+/izWlzPJEteIj0u5rqqH8Z4rfFO89syduy4cA6PooH21/hxOp0VL7yh5L
CeIc6kzVirEzqEzp70UsQz27axxiIP2SohrpcjqV14rP2NpbeJBMJTUrOtGmmyLO
OKX8RtjOsZhTHWjyFgC99RFU7BxGip9/tZQKBiMfp3fQqwFFzrkZl4RRz5v7759v
XJ7rOzTPgM8pDsqgLuI4m8qOgsy31tvD/L6VmsfQR+L4wCAaYsNVyuOM01r/jWH8
bm76hseMGK385Ig1ZKYbz2yd/Kal8iiE9P933RQc+gEuQVAxENcf8tAHRMIUl3nI
k2nt+UvGWEaZtWZv//hLsJ7o3vWFSxVyKi4VEdrVqpd9yGgFcnKAmyd7Ju3MGZMB
DHEpvN61x7bY+inKm41py/h/sgsHRFOTL1zB1OLNIntYrbmDTf3Hhn7E53j6MR+1
Tcf72Im8tf5CzQtLJY2yYHQw/Z7mI91aznJ7BM9cuaZBnVgtkDngrb/X7d4jXWdN
abaUaPrtYOy43QiSP1oPyI0H8Wl5Xr8nGA/ROwAPaG1dvlFiBr3SSAlko9heQLSF
toy8laI3GFpcK7sbePmRUo3G9Z5AJSy22bsPueXx9NFtsnD8GcPVqG9q3Tz8nfmM
lOdlOCL4AQY5SSqonL/fJEKardR9wtWLegUmwJHy2W4SjmpyJ+Lrg9ffl1pFyvNE
Z5EBlMnFzbAPdJSrNHU21DlAcUH9UEU2BAuOnLXuFUmWAKVM3HDtx5EwA8d37vkm
54hzipbPqUdjLZ8Pli8zutvH8V1AtbwAe5UA3aB2BiM4XGh4OC8A4Jfzj+vCfupP
rAp1Aetg2LQC5nnwWGbvA/iHmObFxr2gQum+mcaeHeCZXiOWWqmaHW3NXsOszxYH
oKzdw8rTjU/vMucftVpK6WI1XKpLHyr81tzsGoHl2Od2kTYqXhTJ0PbT6ovGVvkS
PK/XLq61EylZnBWZBlgaWiCXuidCF/VcsEj2c3c7rlw8eK9tAImkRbcftn4OssPV
Pd30dsnhCfStSXAxP9+Y3u8mHECYSDBbDyMoAZWf3/Picf0WPgK50pCXdlijpSsr
bg8Aw9zODZpVnT3lPEyi3DCUPLHdJnviopx1dJSYBIGuc2bACr96rLkaN213BadN
p/5cVPHSABlcGqhN5Y+3fDv2nBqcACAL87XEIeRvubBbcIYGOWja42S6AuuzcK6K
C8HzLQ2yGhpTDQqRhlfZcp7PQrWYUqriIPiYlxVpnGxl74F2pV/u9Uka5S0Iu2DV
liIBXvsqz+wdLSzySBzfSNiYnjPHLz3xmu6izLnfiQVfFyDNQ9HmT6iI9qmUZf+j
wiwwT2BmmrPVt3PTOUhUbw6vsxuyAYUMyeIhr0y+xIM8ulz1oP6KotLkUPUJXYre
jMiz/SNT98nItVWDa6ExuSh90OocbKTQJo8iTh52a4IwfS5R74IKgRARrLBzNKfA
QU57R3J7L6XpPj+ApjiSZOtzHgXzJXX20NfC6CrVwrRU50xyZ4aL20qlgOoyQUhG
MxuEenK6Q2Rp+vbxkGj0wMy8ukKsmNG3cM3DrG30EAy/buifBlEL/6YLEf8Zcmag
hd91T0qgFZVKzGRMP+W1M6npqTvXtWsV3oSjUDi6LXlyySnIJxT18sYra/zlb3YV
ype7c+ZsiS1qfo7677/cg0DKF9DjQHf1Md/tmYSbvht4vAqGwcycEfRlG2uOkoiq
JN4fCmFsSEBZkf4pz7Geqd5/uNg0K/oPvVeFZDnxiX6R+a9nPYRRdsIAhtlpGf4f
n+wdn6+uQtJ7h08QK4puSvAYFu9kjgt+lgvpZSsMyVFwKtqCb5VtOfeRmfjYBlPg
KC/K0G3d3ryuViLKRKTpmF2BY3ay9/XcbWMktqQs1J2Sdavib043d1Z266wYq0oO
7P8cR26BFJf2Ha/l14iF/Oo1ubzAKiVYtaCQRaP5RNn21LN2phsI7AJt/YdsPigS
pJWKNEwHnY7bQ8qw8mQnbFUCLJD5go5C3SMKvP9cZCUDuPTgYjrQd+Vz5nJvr+yu
IbovKU6BUM6BbmzjfXDTychzBQPY4cJE7yp/+SlrtS2rOgzf2LR/KZz5rrycFCsB
NfhAv/BAPFhfrhahoOoLyZP+nTlaCePTGU+gv+7obWiqX5L8cSUSywCZT/2fJI+P
PVUEis0YUIXCN/UyYSMZ8Uls1Nj+3Z6VeH29DQp4w0zfNwS/dzizajNkzabMUekj
mseDU1w7keP7rOBS6kiOhqsULEPGT6PHLn5oh0ohTBluhtLLRiuZY1Ha8VZi3CIe
fyk8vksbdUokSxQsTljVxsi7pmvc935eVouSjZYFlB0LuAO10egAU2gsSp5atL5N
/SmmS9Ly1fZcoslskRldAun6O4lgM6DVq8yF+3CNzSeM9vPU4p0pN5KUz8+2Z9HL
KZMXSbYjfsb2hZ1h5CWJSV2T0PK5l9KFu+6v40BeBOPiNozlO5m/ZxSS53njEmn7
E/vVoP/Qc8N5y330viA8L7ET+zKQqjVqhdJF72CukRmGMpscYo0nW7tlyPdObMeJ
0qyLipAU9/weCZ7BTRvAwvkDuwh4j78CI/B6U7RrHW4DlaW1522cju/cV/C3iP9G
y5VuEYY7KgOEoNfNjXH74pxUR7Cy4x+6TZ9xgFsf8lh8aZV3g+hEv1ORCeVpyHOr
48d/nKAXWbNk3zT2iwY08pZurFoJH6gA6x5h+xkkwnv9Av1DSf7o4uyFlpClbQND
r0jvQQjnHGMgCyoptaVbt1CI3VtUkuStqi7jDcaX3SFOgu//0uSCz820h5TQK8yv
n/ODwwYtXTA+JMTbNh8J6TB10195XD7XLm7Y4jXOv33aPnCv4QsbNQ7XNG+dVb4w
GBh+sgb7it9quLicpfgvh1oH5r52k/9/KEU80thKGtKjDCAzcB+91/LCzZYOpV65
PNulUS+IjFohZtEvQ8nM2zxJ+L7xKKe0/EjlRzVLlr3dCtT5TWLEM55+2o5j/oiI
EXAAdA2EXaqyuaNkOq3JVVYsSWdMgRJupG8Jon4PnvtuTdnXYI2WJj/XCJvVNg4+
7MVEGJYNLNtggNk2T6jnS2hJI3b3YtyIRH/3GFEDNJz77e4ir5FPPKr9sWhvJBH6
7J5c0j5chwgcPCDcnQXGWIJx93LiunLBtt2ndChrcd6WpFKTPLnqNW9+gjHCURsl
CzEDglju7kDRLZ1eJ4K6ztiJI8E19XtQH4O/6rYUaD7ilEtuKLB2iNEtz9KFPSiz
hpiEOpdJGSuKZWBhJSof89EBuE38ApX7d8/oQn+QQI8HGIsdIe/CZTmVI75qtCRM
IfW/TOAcVfXc2rA0RTdBcYRwD5rlvJ/XPYIcTacW0xsq1M2W7eaTGCzIzsUrXaYX
4Y1cl7cFyEso4boiZICy6u4otU0BYPDrynFvVZ2vqNVjTmuHIprhPKNehNSBflpR
jFoswStGE2Q59kp67rSUFTxBQvUPegU9ggzicjnm5P2dGy/XimfvYlKeymAYpHDE
i0Q1ciU6b82TlKBjAE9ady4M8Ogs053h/oAn14KHQHUUzvDWm94Q61dtDhHqFQnp
yyr24iiOXZq0yQEsOdy+eg275GDm8ySr9dUmVdHSRfM1wZhNnr2Z0hjjSWq08e5x
b4RUIbcshoXkNXbWM5LMTLqoZfIpvoO/4QJEkj8q4z1Ttf3SxtAuqEVFi7J5M/Eg
GK3md/ZY//OzkHxBbcFJnPd6z8zAeLdyX6oYrWkVRDQK2KaPVCAghX20PxlujYmb
waACNyCL267apE8NYqM72e7b4ElB2OMSYwExeGWDMwsaj26Ys1+1lXFmwaJ93z2L
uygFuUIYD5UhUfNg1qZOlNfCaT2c9MhYOMP5xSWoo+TylB0XlKvf3nxiNNng4w5b
Mj0CD2dT+GLluMZWjaiRH9SSpky8yyVMf4jLsHTi977pVat2Zu/93+GIgQXQuF38
Z910yfgiVslC/rYwWJuHRBq3nt1DuMQx0jn/10NG0VztBjnslTl2aVioIzxinzjQ
bqQLJdX50nZTop3FNdelAlLKZs5xOR4Qo71wK9gOdUD9pL96ILYKVCL1e9HLlsrI
m/TDvJrxY/PkOpK8+9RmzhSIDoAUzTGdLELZbxvtpTeJ4SCvVxeNYLl+2zR21827
59uKA7+c3FH5g+QSzyKBCm17hYU5laCU/lBcfRekDu71uAjSHnTdpjt/ZEL3NrEN
fAEKKrXgwR8iC3+W7YiTgGDC+wcj/HVvTJMYo7tJvcHzRo1m/oYLnKktDsRRGvW0
oI79rocCqU2f1dhripZzECeltDZ+78WCLwXYjDdwWUejL9XVN8nnBe4ITyo6sVPh
9hMzqNP9ZSlFmZy05NnFf19VwpomzQBwCCQ+LHHtDY7WMMZHUsaBICDXAMt95ywg
/DYKQF2diCze7Bh/oa+kbViUBvusY71lPJx5nhiszakmY5W7I8ErtRBIi6WCiFI3
bMwvGYL214dhb/cm6WAdykWZhEEgNDbBFwD8ljzTu6JaPRP+w56QGble/kZe3V9H
av7KsroaZLnmuYpWWOF53tP4ogFS1ti4RDWMz0no5VVUmQBJUBX3EMEwxlTekQe+
tD+yTa538BMszTzxyYylXMeBqBQfdALG2aWYelrrnFeAn0qym7iYrSzrZ52plRgf
i19CSuMYkersE1S/UMam1zzi3xm2SGOsyhtyZoLJ0/X2QZKQNADzICQtoX+zkwxI
+NeTsv2CZb6ZqENWVXe7LlzF5EMtfXZgCk6pHIf0AcbcFpX2SrzW56Fkuy5eMhHu
wXcJKNdYAYPt7SNyVT0hzvXG8MS6TpJpvLnG4GjNGL0dTZWc+ZPVVeDVhgRdHv64
E+68YywimaEPnHLCV9VXCnoJKhvptL0Mf5Sqq6Zib/rqUqBs/YZoN9WVYFegbfMt
QU7VAZJIwzOf/eLT5fnbuAz6GC1cCQ4NCQKVsjXMsQmi5Qf3cUsr0NslSGVhOVei
W2zY8DBLhO9MUQ/Gw+EsYpl9WHvTMjP60n71IyqqnRWdPhCDizdUPZa4ANwMUzpG
YWOfHEbOlud2ZMY8AFOcytI2yTAzAO3ruNI1xRKBQEYZMULx5VcF2ecezK1nK/xS
xW1Ap06RAhLvCEyuhyLEb1eH7AvRoFpCua/aP0TVrtCoNynEcPgIXYkYBbbNoKeG
B+A5W2yy0JTPaxK5joQbq05I986uHuJ3QZAzLhr7BjVOyIy8BsVA6Ff8FASZAc37
5JnQ9JJCg7aDfMNJc9avvM4r7ZpYaONNcEU5yVvRtECyHn6iteuPm23FICq/Hwdd
0xW/3YtrJoiyaIuMuKJ24d5QCF73nz6ZzReyzPNtBz50bthjhrFYZkMdFgyxxZBp
oKborO3WyzJJfVXLP1RgWKyNRt5WybB6n4slCt07c+21Sra+5SXhZnltwxQeVzZ4
3NvRlSACzNrgtuhK+8X3ucrfeG3RZoXXyORMOBwsTTjpipM5EQsv49eFwRDT5hsL
RndrxveV3K8zyOtbSId/WgZABeF9J91L6syzI7zP+srSVV1VhH1ZV87qB6S7zTM0
3ls/WIqr0WzfhohyiU8niwV1tPBa91MZCEkXb0eOnJ7RrNpideswzGVSzq2fvYme
EGkioqCox1JPZMCjtizeGkCNAFBNFxei6Fz9EO1U8aeGFcN+O4zeY8hOpjCNTTVv
mVQYaCLEw3az2GcVzjbPVBfXR92nisUZbHyYL1gOTv2caMcI0oWfuShph34lIyHs
JNyzrEVUr5/mP8Zn7BgwnaOf5ae6dlx2P5mJLzxny8mG6EFTLgjdgW/5hSUEj5hB
g0M1pVuDddH+FTCjC9NriKFywwoU8hjm5RfKUtK30zm+x+knMc7WgMkYTXkuccO4
32z+BWx3JmuKGbJSAvyVJmkj8n9qQhSsiM0LDrotr6gSdofsxVDLqP4+//ODWlJt
Tf6XhEb4bw9j9VsZvos9ZrJecWW3UdTxPLb55MsRwP6c61UXksMP91Kzh/GKmfeX
Qtua5Bk+goh0SlmaOwWNUUB6n2F6THQTab8HR3c9PWfuDrscNwlccZ60ctBtHAz3
sb32d6ZVzTFARMSjxbOQbGOwvm8vd4WXv3aPPF5BBwuF31lnd2kz/guuISbB4wmy
Ayadpl3eH3OBKboV19G6ysd1Mn+IokrKPWcB+gM1pGDgBmLgXOZsqrx361hBGfVQ
ARSCjycMwsE+4D6RjPDcfwlV/ZYeIkAxHBRZwCuC7BMHuaGHICFMMqxGJHpl9nG0
LKDd25oSpgjo28oWgK0Ph52hvlYnvhlvt89ZESaB21yzjlXbf5L8Qe6ACPLP1peb
MXI3lKzR1pX0oUHvRYgkk5sLjWWK7GTv0Jdp+53AA0eDOj2wO5iQXu/5C3Djq/G1
msXpOgE8cKwqNOqKXHNNZYVNtC/N91t9VDUitSSbQUctOzzWGFdPT7SzIX9m6VQi
MNtNkA2KaxezGQaW+vUz49PIfLuib+cMNIrQ16s/8OxBUNl3uAJntoRneCG1OnmO
PK/CrY6kxxJzP/ei45n57dHyv90xUb5VqB2bqMpnklWnOTPne3NfSJGVV7yqeWt4
HKIpnpEEwyqdCFrlBpxChrU4/sNwoILfLr52CLHfwz4eD11/nx1YXHBs0fHHNbv9
6AfFdvED2EtXzxCcJ/FRU/3+ihbyZBBPuRc/15Dh7QA0BzK1ozoE+zuUDszEhCF1
6/D2HjgfCteQ7jTIQ5O1beKJC+dhH3qNUzRnGz93HZfkBs2hyGD4Z54FjKv/1rom
p8RUE96L39UP8RD6L3bwDMY1Kkp+BXO5Rv975F6YUBZ7yZ/YPXTLXBtLrZx7nDcK
E8oVtldppi6NGgejOM6E14yhAjMQoSRyhsrOLsH7m4NYuU7KUM5/tL0cXRskVirH
OOCfrE+kfQQPFpvH1CgP09hFX/gY0lPSblky9GOT1pWoqSG0VDKKaZS9RJ8Feskc
CqBS+uaxI3atXrLoIcztqNlNIrfnQD+Lvyg4FkcDggzB4TOC+jpwzePa6NeUV0Ms
szcnNDsXsgmISULIFFzlzY9ympA4iEwSpe+TXBRN7AUJrYguVGO55JuYCq4vl/Ju
h33VJ0tUUSAdcAa5Gmt8W/gkmOmHIb35cj+0dbArBQXxGQhyF9D1Seulvk6bXyts
mqJ2vHnAfPyzZ2StBFaqv0d0g+snFBHOhtVYADAZMCrOGrx3l2K+Bhu/EILhNuko
7NnuhAkzvrEFGcAO0S/BZp7Jv3Neb7eSlm9cTGtQKW/WJrfAbzt3CCVyZq9No7zE
rV4fYcQTBIqv1C+mNjxcOz6srYrs/Rh38013bTi7mer2jD6R0P4YM1ynzLUo2JWA
tHcoT8BcSmfXNPEqZEYPMUtix4QOry8J1x1+t94kIol6vlu8pmrVm/B0l9XOui9W
rmnBUlcBLJ9IT8lUG4kjiexYZRpyLOIsNYxaTw3+IE9A1nAX6adUi4Is2RHybrY0
Byf0rb6d4PYKQBGSeH9omyiu2+4hFNFFh4TherRdWwKcDB0PwcIQ6gk54zIzt6U2
bvpWUhmTXfYhI4lbjlbg7Q+fpil+0ACoZPT38wqO/DpXM20FGM1P5aL3UVqHIe3k
QJ+BWtgfboCQ3jGKw9tQbz4yOEsg0J6Sb4oEVfvzrYbZET48wfZ1Ma1DAlZa2hSD
y5LwCzC1Iw1p/2T7LDr8xpSf1n5y+4Q6kPFdEzKzP+xuZVpcKCffkxKF6PVdKtbs
Bxb3Em9Ev7vwVcNbmnwfx3q7ALObXzsSkdj0UVi7/SdO/JKOP8fhaKSHn4soO6AX
ZXQPpKOCT5LGzcBNVdiWt1j4rhLy2ka4P2R/cb1DSD02lk3p0EWNhzljHd1otEnb
abw9H/JpQr1Qctb2GiXrNtTgkmcV9zxl0dnrXr1yXq7HPSQQ2dXT5KIXjJHwDVXW
JT8iyJSbMWmOSaY2kHzYbMLemf6vFcRkKlu+7H1IBHSZBeKsJ6NWg6BiNCch8lyR
0JUUQEJ5KS0l9QR6/l59o6GdVSPAOD9hoYlCuA4kgUXeedU6aIH75Kp0IU+2UDwA
VoC6EDpdr6ciDwKJFHFi5WBpbMmVR3qE87Ce9yaDZnHopQ0PC4M1QwvWlH6o1s3L
BOUg5zVA0UFxkqY7jVaV1OM2LJG8QrSYyaFczdlG/gopn30HewbCi2sdkPPjzmJx
6RRx7gWABopr+TJUkZcs+UhJu3ccn/d4N3640xADn3pbBWTwG4Ds4iyvmogejC3k
UJpQndo3+KTf3Uca89o/novnXWhOlyRkhqkvBq+bFrqRu5g9rFZoXmgTEn+16u+P
1GCh0BqP5eiwcWm0703UrRuojEWJ5uUZAMoXe7kDoWuRL64J/s08sJir/cRXeCmv
p2HkRaic8iDIw67ev58+kKLZX0/fhJAMGemqgUkSujLfWm7ud+y8PGZ8RwcP1sxX
TVuCIcgelrZz+avHYmnXBNiv88I0IEaDblGAhO1Y8qqFVIqIB9jJ59K+Cr+Z00Tt
fH2CNyZpJKvoTilvpT/2epUXgz3rIKpj0jckJxCLO6S3NhQhCfRCgMsslviyCxNE
CC1b0NZnRj/sfKTpWAE4z0sgQ9lIA9EeosAl8ctic9WBXp+BQyYmsX6TKW0H1Ojw
DVuHK4YrF/73bHJpU6QWp4mvw0Jiv/wtGZ4zSP5g13YBBTsQNqnJaXNWEsDiLEmL
4uP6JyaTfg8DN+AOP6OufOjh1F7Brs5kuiTOdiIaK+3KbaaXNerH5PbCdVlrQssm
yIG9W1VGLrG1QxehW2R6ASdR8JRsC1zDOLeCFAZy6YqR2r12QylbQNmrvQmyo9WI
//0CQMUe0nJZ3GI8af7YP/8WKLSDPgh01KGFdGcQ5M/bSJZ3JE9JDGSgvl5XC425
4BqQP2NGzZTDz2SpLiSinPDe9HKztWFTQof62vXV3wvMPMqyOZd5j2NE7ISDhvfF
FhBqdnc6O3IEZApKEbdBaId5eHqct4y04r5L19L8NaQjwYxTzzqQvyGUEIpo7wLn
Vccf7Nn3Hpns2I9AoFz6ppOq7xgTSDg2/5zJ9kkPVJ0JH2F1VPoUzUHBRP7O1yhx
tCh78/CBJ3Ktc91W4jximpSjtwn0OlBusIS0tC5VuR2yC2QMNKLPk03LPO5k3dMn
jo6ts8RX2HR+rOECLVzxHkBbHspb9DlKVAIegzpe9y8uTyT7udofBARcXscKV3ob
EnZy4DSpyC24yrNNki/IyZBAQaEf4D1VfCytjeXpJdyMMVpMH0DqcsNGUVBEILHh
uPSk+2xtZUQwM05kFjcnErNdq1g8vKrhgFKwPW6WCEdJATIhzvzLhEfBHTsHmRyV
nBS4nBj2jfUimblHyxr+zvCodT9i8E0HlJTYKEhZ6OLJW0twmfJcPDSki8xCE7zk
q/sAoCFai7+P/2IQmHskqQPCLIw0bavBAUcfaG+ow5zB0eIMILjKNuyBYUb+Up/q
A5AEEutaKBN8lLNcrHEhHnOGUjbMzTGBaT3WzF6VXnwq0yV4C3dnFg9ps1N9eCIw
gQQWxYwoo2ylXSdN0PoZ2vLAhqfYiqyb31PC1XykWH6t4Zc43NAK+iog4WNKJr3/
8bl20S9dYpeXtHaWhmpFUNzuJf2wf/RJS/vF9uC0AfJXvv6ApzVFHXhBHigJDROw
xlPNPrqjA8+K0A5ofpOUYtyceWLm1gKdOi7ket7KDoOV6YkooQtsUoZiLaKTEpSS
QoJQ98XR23Q8XLmGjnx4m/qvpy45ftz5Z81XcYTx/Gk46eLWUyflhVNIV76DMwUt
ObGoOx2W1e5nE2YARAawi5/XIilw4nIXFmx4QACcrLZU69D7fvjV0kkYGuv8KQ9J
eDog5LSSFHnQyt2+Hzo3tH+R3ycMAb2pvfA/77pE5Qdq2MNq5T0MB2NDKgnLQ5er
ExjxrQbtQxnTJExrr5hvFlhGT0WuvsnOEPOMf8QMZLCf5EHMvp2HSCIcNAVLtRMZ
/UpUWfMquwQoVE+oeWi6W9K/H0lBNLF7xaaGZo+M+rx/tnQghnnzs4v8Pxd+RBNZ
gyJFZkn++MgGQCZdzqn94eiEYM99HD4tU/EmNRqQtqVbxZyD9jwrZQReogB5LvPr
FVH4GnJTaykExtBaRe/nFEN9b3OwKBZMPpUPes43HfEeTZt7IsVoI8hiOLDCm28m
DY6AyTUJMY7GRT77nMWGjKvqlNSJNqAnfCl4LiITMq6PwK4kZeBKos/GEtvh/gfo
U6Hpjv5cnGw5tKnBOV2JyE4Xz9ow4Ibzng3XD9aEdldIFt/TGzLflgdrD3KHgdFE
4IypfvOCKrOFUq+5tNAfkp2nlKmBn2aGqYzOrW1na2S8kUODA8jz0X3f3zqh21gE
VtYA0UVcettnU6ievgttlR2ygo2M8NkTn/bWaqrmzJZ22zXObZbS2XnuF2ANwo1+
7mtEHRJHxTMP6hJZfQCCmq0y6qS44sXHeWq4O8Il8pqcap7arl73adgqONxT3Kql
PloUMEzH14vegU0jVvhuc6r87xGs6ULwutE1wsfo/iRul6JorXEvgSfHWC+9vfP9
kW+xmdnGYIQsrS3iP7eSRNp0sH/IjYTLsGWV1219WRVpMOHZwaOJOVCF5kbWdopq
6Lxbfg0aRE/+/lYPURycyx3gmSAeCe9D2bLDPVL/4pRtjYi/14AXMwvOan7AmrEK
2q01hmOdhwmpBUo456yZGO0wByGPDAToQTcD29Vc/CehSjfP4+PsOUaNOUruiFUH
8hntZrSsL/sEWwU6fYHhISza6Y2MKNrhtfyzY1V61XdeGp+28N1W8r1XKXYzeVJ0
SHdjvPKXMgBQJwziSOlNfNgM2yO0RPFvlMy+EO9yTUoLLNocLUyPEmjJ9ig/Rfjb
1aDJGd6I7C8ysNjwFn6qNwUoJ02B60uY4LTJn/RuEOWHcf0WaJK+3PlEnkn0F3Rd
tPDizXJ5qwqEJeR231IwHrNwVh0PTmrg4aOt+kdXpTBQB9qup5cP1/aCsMOe9WYV
h/+vGQ3wCpWMRv2etymwJe9peLCJ+e+t0/AsbRulRnkNNjo2XwUhSHGGHrplwYVM
4snyy4F9DX9UJ9PXLmGOEHKNCkcCEe3sDjD2EYkn/ZIrJGewiajTWV+n6afsysoy
jCf19562bqugs0RJBTtd8YBhmCSCu0ir+sMZHgD6OFzDkSOhCgFLt9kAMbjafgm2
9f4+OCE7KNnwupGjMmNs8yzpABT0EDgXVQ2QQB//ZiOkLWVFXREsDqPaJKQqjEhh
6/73sTLBligLb+ymt2zeuATlMIXdaciNj/lG0YB39v8kmpX3VhLnu8u0bu2fWJVW
+BJKC+o/8kY4VRQk9kx4ZS87Wk+OWAPfoqghXc0xViCpk7rz7VpyneVNcPqht/Nc
cRIA2L9xSTSCVKz8EquPW+sKYLiq+pb7iOxo2hZrBi8VoNARKYGojNbxOb0d4x+j
1mP8DWiC+VQGDwRl+N6jNHAq7LIWWRODYFWuCfmJKU4ajle190/9gxeYidQjFVNc
r7WJ60FtZGQUglBbWhKgz0s+AQYE7FmCKInDyBgR6nPZAyHxmjGEBV0RoRFAi/Ps
WvfvU7UD2+I1y0S4XDYHDjOq2sVmV8mvf9W05zq+HiaF60stWnAkEYhuA5gSzXDV
fRvpGv2l1IWNMG69OkneNKQzofSCCmhivfMd1iuajLoJ/aft9dnH/xKXUA8E18kS
oo+QYmSYgH+kHvo7Km28qKH6Un2UwHIB37HWR78WjTNc0H0Ef6UGjFyt+ObqBa9g
Gl/CSv1EcetT1a9+GxoMJ9R0y0uY/ON2D4trO2HjsIOVt62o7B8kNvShpuuuHwVh
CJ/MZEXMonGr/6UNvt478QGu+qtJ8KLUEX/ew+Lc1QtbABgkCJAH0gAvzSL3Saeo
u+otgTeN2Tv7wV/3cLqSCQ7r8P6km5Y3iRTmNQ4VTyzzlj5tWxcrOL3QZS1NU005
PnR6kTNqIy+5lDjjAlUw83edwgbTY4uX2P/HdeZ/Bie0G+cI1RMUHBWew8p0ybDH
ctlPThk9p0VAeKSqwDc3dtrFvTG1Q5Q8nLrnBRm/bQcwXnrWpMUsczvwBTR/mJ9R
pyx3GD2u72UY49dY6NTBCZ8Y7SeXncEFiHAVmMxirZLlJGTjh1pGe04+n2VHi2SN
JRBPZMgz17Iz+zYE+hsO6pNu4UAyDnFn2ujiNxfcSQvivpPSRI009nEFHEfNx9a6
v3hOQpHbrezq/tmrTmIdFsfs359ZKBWuSvofyHTrAll+Z7D1qSEVNLRA8wgOoPmB
d3B1e2q2ciT8i5hl8I5AtlLPfWem39QjHoxn1v9vO38GrjgnLFc+OaGnJHBOiOW5
uofrc7QefzijiqGBQgqf1RESD4z6RETbYmxKpQApnHYcjcYR36hBOMOPvuBgyt0+
PLDublZLUkvZMPBCepK/4oAUyL6UqNj3CKHabKnAXOqeJw5lI5wjxCD43pQa97Nw
Q+6GD7p91v53/ZWZWvb/ibZ2BSXRnUq7wvlyPbtDB3mFttWCO/FVAI6htIiiE/8g
9WZ+xB1zmEO+iCwJSOYsVFX5PxXh9Ot2LjLpvBOhdyxlOxg+srDzVWalFC2TBta3
ajLnszHBSVGQ1uX8scQKK1kygw4VduvjZbC1RIydfvIOD4PwPhCF8YhebLuN02To
6U5LhlOj0haluzAvQamGEAXR1wNEeErZK4QgYA/GzwnB7dYLThnPBhI0sj6gFPgy
gTH8LBHLxk/O9N52lGIQMdsE/PuP6yDDOFt2yZ9OyPfIhmx4BoHsbl+iKij1b3Yc
Ff3kBslmovDlG7PJmF3yA2pwtTN3VKN7H5lFpVDASSa9q/ISlLSdF6Fc10UR82g5
fA6Zn6O0LM+QouKc8KQJqRGrvway2g+js1QUenGZepNTc1kVnL8wDPUFBhHWB2ye
bAelnlReWcxCST0p+/Fpt8jbunlUD28vpF3EcDXNJfXbmngNKcKbao6CjiCENIHS
imeEAQmavhcaWO247FnDpCKsRhjmepVL3LKUPWcBNxUyCLkUoK8E6GNg0F5/hO8J
ENx/n9/aUNjmIU7qTg7Yv+JbH5eg9zokHVQ2glhqmg+EMRG7GZJ//nLDayWro/oT
iPzw3qQHLwqMa5+okbYiZWDFfU8VeamYmK2zyxS7AjACDGk86z59W1v/MktHn2Mv
gbNCkOxUynjNDuEFGVnDJX90c4/WywvIZRSIcu7heX/feK9FREB9z6IPY4CvTiZB
5x3TVXyl7EggS2JLo8PRg9ALy6AqokMG3XLXxqLTeGADAusczDfQYfKIjZ3f77uc
wdD16LVF204Ih1weFpOG5EjLVOxEbNbMwh8kH+duaFe5Q9FMA6gIpZd2GtXZbQWU
G/RDHtCU1L4UKpx2bs7TcdJwc5bWp2+YQc0YyKLy5cICp7z+uiUpGafsiAi81aB/
rAN8D+qmf9As1XGbjd44tZfrActBGAa+Kapf9tTaxbh6K7lCmD1SR9vChWGCfbJn
iMcD+bU6skJ3EQiwOPMyYzPheoiqNOBsPJ3IyPw/bQ5DiYRl4bs4Vh38VU2SssaL
dau2rj+KZvUI5aPZjjINQJ/g9k7PmamVZMgY3XpVharXA6e6pKR0tMbnm9UcadBf
54ZdBlozaweDBK3CMuXhXwfCirsPBOioOv071LJRWFwB+Cd3GiplG8LrfNuNxIh3
TPVFPvwWO5C8s+17ItGxnMGkBtlW9gak6hpSQfsWzt9XMT67xNHzu7zbTTUB0HaZ
fh3bFajtwGD3UpFiURcK6DxPm3qFxZrpXmgEl0DU/T4GhwJWdgBa5HXsahaCkmW2
vlj+WB5k3xexbIxdKJ37FdO3UWTEQSO+QNrvuKOZLkBc95+HooqP/VDNJ4gbNej8
xY4GZ/FeMQCMANG4oOsvHMnkKeswyiwU3vsB9g6MEgp4G5rx0qtFbJju+SSBGjik
7uUmHZGA76YWzmvQzxtBTJZxRNb8iNsJRwu3XwEy4jB0tuOA+z0VFs/4w94410au
korxqdbKnd99wnBeqSF4cDrAnRTeAwV7eAqTtyKGd5yyJqJIQBE7VDs7v79Wp+rK
IaKXkK+y5PkCs5XMVHji/Y3+t/FixRMndLDpd3bG6wAiC55XxgSWvg3mNMqZ1hzN
jAFH+nTvwldLlWyzlRmvOIfE9X8kW9LlFztsvAe1TRFCOT8YxM4sJYvSgYnSKnZz
MPT471HgEZKLTd4mCXibNTGbOWyatt3sOkMoF8tN5SR1bt9ciH4ZtgKdLfINHB7Z
iMio8oSpZaN7QZrljOHTmZrPFP5EeoPrHmMs/++j+OhzwPfQnpYHDgi7iLMoLLSY
EzQUNL1sri+3f5PRnCcZMCFbAHL4o8FbIaEb21IVpOXT8Rfe5jrTw1vgpGFVWW9Y
YFPQg8SntUVLF3RZVC7QUbTUDHXsdFoXqca900ypKpvu0NZ2ykXTd9heZbRCtAzp
3vHLmsUs43eXVLOsVBBMC0LgXI9QMeEd6uvqzpyuphbiyvskkLLDu0ygd+tUchPk
oAwrijgdXDA79nvEz/Qm6xgTp/5m5G41EXPhQpniQqHyKeOE6dJ4y6/xD0f5yRUN
W2jYEtb/e5TEXiCIZEResYo9r0hiX35TktKwEwvWxAURpjCghHZsIPUBTSjrilxh
Ya5Krpknbr1kiNUho/y+Aprfk6c1L/U9X0twtJ20AD1RH5dKs5SQpDcpYZygbYAQ
nLNhnMN5rOJi4aXIDgl7wVNpzsV+xfACzeZp/xJSndxh0qDBWCd8OSbOcW53FBIn
iqF4pDY464PsO99sQSAZ1B7MMAkcTzmEbsMg+BM4ssoGzmq/qFV+XcKbgfLjgUYO
kgzpFkUWcTYxibTkEMo3yyKQq+ttwwQMqIW9SE8oj4815cDGlXk33RXmUs3r+hft
k1L179QUspFSaEFLlqbx/bBDMarrHQOYIADzdS5OWqF4kbRWJitVyjR1YmEWQal4
O151xYnuEqeCqOTkDL3oXbVStanCMs5N5IVi9Wv7+QLHtZ9cvecpaezUuaerVSK2
bp4wK4OhEHPaM+CTUeR6FuBa1Axh3iiloUrjVnyD8sj1UmuaOVQ41DKd0SD9ZcFL
HUo6YPayzIiCwUSxAcPZF3q8NAE8CGq3eXhkxUE7b4+AmQc8rFq/7bEs4Fip53sA
fqBQqkcLrWbQq+fVzKzlK4whG8It4HOtgJUm5woLRYKqyYh4MVetORnk7hWiQ22/
Zj0fW/DjxWvZa5PDdfS6O2eKyCe60LN567gl5onxELw4gpixthku/TFa9EmIGDfR
5FBRaKHBbWonYYVlIGaC/QkIGe7OuGzIfxLDxG04YTdCqHc612hMfb6YSZuo8mdF
e1Jn4fhJ6UL15z4/nhcjZVv5CtG8rQvMhl8UarDD69bB7MtjCPCTl68bXUkZAoyZ
F6DeRcITfdgX+V2gVzElRbOF6fCmFR0UpWHS9AL+6d6OPJjQ+8V+IcwPq1xz2REc
7SrL9SiVt8iXulPYlixdCLFxdGNEOs+ln8PaIsLeaCSVQHn8sjTReYXZX1cXtxJ2
myfqkwdjEUJzrULYTPXyRaJvyNk0BrbknPgnp3cNSieGYskZ+Ez/iHRkUvRUvOv0
z0Xp1zDgeWpM08s8Cuh3yfKEi65aM3FR23PfeFkJEbdV4rsrYHOqKDN0PnGrfE2R
HJFVFsmXyMTJPMiEDtxjoU/y3vBCoxkrcvm/899B7RIbsUcG6kCtbHbQXjhyEcpI
XrcXzk8nLvCczL3zgfGcrWULCZVH9u775428VpP2uDlf6pLp5HIS4Pw2ft9y9XtF
n4bOzQWulhuOQG0bKUl1GjDD7GE8vLdO3S2jFXV5+GNeK39F2MR4t4ffDTXuHb5A
+ouL5ajcf0iTSplR848gF8I6Sdg+34yU4JiKkNcwAhn4GjbYR2pkwmXD47NzLuRg
lauwOMDH4aC3eElNi1fEaVMkonYB7M4KHE9SjmZuOdayeXoGIzT4PE9JqtVck34L
LpjT1zSQGB7qsvB0pY7FGDkUjduxrXBDImRkipGJx6JUOUW22kOOTGkB6JyYfNS9
cfDGjyj7MSqdxWjq8bA0pCRG1ONGNXoBzg1CDGf6bKeU38gsQJgsRzJ0bVQZ24uR
ZHOxUzk2u/nmbMaNbS+zJDdQudAq5HVnuf2XtV/zCCDCZXQHrnmUcbdsjWjZB2fo
SEKgrvWfF+0GQpBxcSd3byclM5pXnA1QYHo2GgoTArK+kjAimQDf6vslTP8RHkUy
3+fgfR5cjLT+pwfFj2sYjXox6FswNHj1NO3OMH3tzpCqxa3oXm+pFgpDLM8V3tkh
ump9PQYL7JQV4vdx9lTgI8uqSOvqb8iwf7Wnn7CIndNE0zrjNNubr5hvHP/pePzt
6UNPwe1Mq7FuslHHkazacLXlGZ3TJl1zYrQqbD4KQKK7S9DzXj9VbDxwlFEG5/25
qFuh2WvPdln8SjXS8PB17J3ssMTaPnYA2nuDmoorvBIcgHGeFvqqOFD0wcMj4o7y
xcZnOoNCMzRXZ0SENzpAZEAN/EKtiJCtkSCNDDO+2PcQtEIvktWhnJ3h2y4Sqqop
11mWlPrg5At0Dt0nDafaDXt33Xy3FZ3lQLGslLWfxwMQaerJMDRsGc6Vdm466kEA
jGIzssPfWvgwbcAu+maQSdMjtNpWeA6BtPS+HQ5Z02TxFfU0mXE5J2J1dO4Y/ZhW
692JBM6tice1vILtX0TGF5BKiB34ewaESfVAfAetQB2NdBAC1vdLJYYzPcsZMzqv
AD3WNkQFNn5eGhYqIWZOC/ZULjNsXNo58jOylv2MyCkfEeRZhKQBpmYlyMQkG30s
rZBQiQIghxkFgciVMJXhQOUh4BMrrdHGSwQ0NbF9UB7f0KKmi0UU6pqo42O5xkdR
dSStIX5PiZUGOdhvSIh1MvChVSbpXW/Oj9IoagGkvWEvujEyUFqlqJairuoSQCtW
yxe6LBbKN+G21tC2gZVHUFNxWcb8GtN5yvY1UfzPczfEpDiKpsbocDNqtgYMTDzK
DTI5lKpEs9MmSN72Djbu1Sr2UZgjZ7gJEX2mkN2+JKHDwozruIQ2ZVGF/1fE1HPE
fFYIKK8Ox02micnXKqxoIr6sqUREHPmatoT/RCOcN2oCznUntp//I7SiC+COfpFj
T5z2IZWQi7QnN5fNq42hpEbxQeiP8dxRLpX09QWf+il7OXFQ2HlM4+GM6m6/uFoS
En2ycN4jlKmNxmzy3cSFR9DN9DZRo4O2uojsLsLO4//hYkAtCGDqO878TmDZ9Tg3
hObNwmybIb4WHm4N0ls/IxBXIz+ZLFErxLTLfk/YHQY6CBQA7d0wSKlIl1ZGbv3c
GzLuGfo8sxM1zoGMyuJ16RYrZJWMQnzjlD2CDaIuINfKPGTLF2LuNo1/6rGA5514
ZvIkpUHDQM3rQvi1XIN8GeohGL0RPRxrot/FL+rdXwAQ9GNB7QKjF2FyG5/ZyFbf
PX3ku32Oc3WZJY7fKp9APpLAkQa3qwxw/Bym2hQrUTuULqVSKs9V+pGAvkqh5mHe
L35DPY2xmVs1tG4JX046zAZ3hUXxUiL/2pqBrGnsXEnf2dBFijA/sp9hxpAUS3q1
jPMT0ydLQIrCNQmz802JZ1Dz8HTN+ImO8T09dQJa0SkygjDVGLm+RI5+xoaIJ01L
l0eSeJjjximk5aqWegrjOfM3kibGK1qDdUzJVMD7r/29easYs4t06+84+ssV28uY
0VCn6R2duQ2pAUvBk15QPbC1p4HPDO0BgYREmdcAQZs/3P75X3HWMyBIl/2s6gIw
uR+La1cH0GRh3MM66/sGnWz3kHQGe3gLpwP8GNuNfPtO0QeFCexX9V7jB99uJCiH
cmA2/R/eIKuBRx8fvPHkHKhbBz5EjAH06GjVZEml1YVS5rISHvJgD9CbnD+W7Tb7
y8lBF9XVmyX1GNsKv7WWs//jwZK6MpSHUweOCAXlWRphcQyZjvq7XO3mXjYnhVUD
oayDKcR4/PhEJ5XPgkbQ365HVLQciiEsJI6IKOsz4KcTJyr2k5hjOdoFttLXmjAb
N9KnwcVp7AyAPJDhSB8l/ISGhUyaIHMxgukr4s5DMm8kz6XKQklYolH9Y63xwrfm
CQbS5SdyKILURiXS6+eveg87TZmkI9Z+ZzJvbXKt9wNP9qS9ceTswk3d2xQ6U7/6
GCSJsDK/S5gM5SUaUJt5MQL0gRVBSZma5Z0hj1TftzI72Ei0WtxblKltcAutoIOa
CyEQk5ev/zdeyCv/jChTvVmHG8CUEKqIeGRDlCTYjK9PsrohgIBOO3QUupTIMo9d
HF0zN/cpRL+aoTf7EKIdTLBKEqF6/y/zolROwXHyYZ7NiqYQKIAi5ItM4DP20awM
5gjKuyru8z2wFHbnurCS/qiXwW2xMjyRQAj5NkIpHoy2MD+FcDTzOCtf6oyLEArP
3LlfbpwUkoYLXDfbyU1HrtX2Vx55Uf1R1uQ2cE+/45lUpxfbRIuMunDU5tD52Lo2
9XFg1sqIB4xnFnBM4WI9HmMODnmChj5uAaH58WFtS9oGAZ9/gQd1WgC5AqCVduCZ
jlSMRb3pZm8F42ooQCs5se0SPfKdg1fjhf4yYSDtwDvo5u8ZwOYRQZH5cSb1XyrR
MLZFNCEppfc0VE8o/o9nrWsgcAWM0k5KoMvZKwZdS3PrZQMKOVXjHcihseN4T4K4
2nS+L/SZHm16MQglS4lFRbCISQ6KVsJAQ0T8AX3wvoXE4cbI4RaRkqIzI4AT/gBN
6QBpaU9EwJ8XGaIT+z0p/USRTS2DOsMd2WKi6u7+rK+FJRMhotLjF3W+KmXR0bhh
ohUOAQM2DEI2s3btZXszANqQUtVOVypKxTsYDSaqcwYDrllBpbMAgATnnwQdB6o6
5fSe0R8Nk/A+uVVi5Z72rqFffOkC6OxlLsMBUzonZ4lQghU4C4ynsYYvq7B9vwE3
NCNb/jxYaoGCB1KPaAUTdjEslWVwAtHTyVza2A7Y1dgSGFdGhNIsia7mc7pAWwk+
zun32RuOSHdELXskceE8C/RU53EsGc97u+1ynI07sdrxZAPsGI9T++6FCIVEDoH0
k9WxloLTwnjhmamTRi+lo5/aQxuFFzpVYFWgW8efaaX+NtKW6pCHtpNjN6+ewOLu
MsTgY6PXOR9Ft7YMGt7HO57cEBvC1EYJRHdppizlQQzeUij2XKIR3sCoYkiHg1pF
99TvmmfjqAMMuEchppsJ5/HgTVTh1SsaudBEOGCYC8ULSJw1WHyK8l8C7mhsp8Mi
vJ1hJ4pgr81cSU60qc1b5swQzgm3q7xa6FiVLRj7hVPoObnpkq0H8AWOs0M6Hr0z
jXM4OFXxQ12dPEYTXxHch4tFUlX40R1G/PluQPBb0SB1QJWXquL23MsZWQ159Zx3
csTLwWuPdshzYbVOJkhN0nSKtuc+SnkbeJeO7JV4s1hyKDGM1U3xw2uY8J33SqhW
j+3trarExdOJIRNcuvM4DZ/9iIht6CWAnwKqU3W1SNzMquEkpQMRlH2hhUEFbeL8
olj5Dd+ZlAJTRSfQwenRmTjK3rmgf+9WdUusIPnhsLrSmAOmiclupdz3Ph2tG7K7
O4fT0DWsvjtREd7RJA440gQ2AER7SnAHSMjwLRcRP8sPT3yadOCxUl/FrnFwTaPW
RyTarqgkCG2pdUmaXpWmkHcwUqD6WjDUuSbX6RfDGjsWj/PQAjr29jeSXzeRRUQU
ZokySqDw+G2QhTEGWF0vLZ1QXEcrnKbxfqvSfC0A663yHG6vXCBrFeAG1cWG2v6S
OBn8k/Actn40yFDMfNzlCRwCIO/Fq0LDLlibIAuLH7WXHzu6MU4gTox3ASY6gSOW
5Tq1j30ptPq6riZAIXvey/Y2pVP8G5e+/PaSe+6mg1Z6rM02uhtvTYSTbDz0iN/5
gbcyOMtx8CvMME4tEPqcq3qv7l5XyhB96VgXU4wAn347ztndyYZccjNS1kIjNMZA
M7c0/23lxZOzBnhBV1cK23FHUjHhnQA8TwKp2QxduTx4qmVxdEGyCKiSZECzt5DA
qtJh6YU7lIHmZDx+pZyXv0U9bThOS9vDmAe6LSHbKvdgA02v1y+GoJYUySXc0ein
l11eCZHxVQU7Clbj5iNV2lNfC2gol8tBb7QNgI2zWu22SmEP2e3d2LZryd5vlClN
KspgCq70IylF7oDxDtrP5Ca7mY8fOnzAmLlshcpkkRBKxnaY4GnFYbujDXhQ+wuM
MQI5BnZwfj/skjMZ8IO985SEzoJraUEgFRmrNyRUnz8vkh8GH3NpnDiuLucDoDCp
SjJNF1YMRqS9rEQNH+i5i1StkQmhPvsTPqZkyXz5KU5hpedpAY+awxC0HSlKXnq8
4aHkO0uUbzz+Q20eLWGdgZ3eVWEzHnVxvCo/DP9F6CrYjH6dKJ9OhBmC8geEwU03
P5AM45JN4PFfFPvZp5aMKosUpzRnBq5OOpJkXjB+1ir40Sx4/h0cSjO8NU9sNfrG
Di+hanJxTlvYe3UldsA1ZMCVPLGSkTCX+7ekkhDEkG8qj4bx3Ka5RsiVLZfFzyTS
2G/j2/s48UPsCaAmHHw+rHq1zeKEZkAbquJFuLfD9smW3/21pCw/6z9of2i8MZrv
d8S41jtQEpH12YZyTxa4Jyr7un0oOhnbzk+JNk0/AbJb0Mi9vaZQYRv95Cn6MBMK
cVnvZbTSiBy8AaOBdOM84gt7uSe6/iOF2V5BpbucUlhbKm4rozL3CC9ff8Si9mM7
32M0XJuwLiMiz7NNjOlm7lq9/1xNPquwT1Ut/mHurBYF/8HddYqsdFDvSugQymJg
8vzpTek0WC/xG25Ra9LBZeRDoSBSDwdMaAMiTCIDXYGsimxfwwCDOYwYldrUFi1D
8hcEDStHSJPXxcxYsrbkMgwY4Cb/VfEbiuR9WwjWp7/w6pZvxWgE0RZB3jAPIwuL
hHc5ZTBWGrIrQzJCBmw2/RiDYvvtdVaOzCJll0+LgaGjvU464nYfnlIc0hR7KMmp
diE0fFYoBonWxxbNNia9hfeDBfaoo01AXgmR5raiDEtlPDNraze8PqX5WU5Ys8Qv
CcYP3277vRdBEHbz89eTazg1rplRL94zSeLIXRzNE3BMT97ph1THFq1yLP1vbr4b
6ve6rhbdMsPWLp096SSB8shS5qbHF7gKXdSq9PHi/yv3r6DTJXATjprYKrEDUAx7
NfgVNGIFvsIqM01VRc3pm1NWA8o9jtLHAFR9YUDSgU0F0moRJLp5wAW/fJgWKfLL
95WkWgO1RrKvBGTER3WTH0jJrXA22dA+5/pj6ZxeqNQWTsN50PGzGtBFz0irH8EC
r08j7wVp0F7dprBT6jofCmoh6bINWRj0gb7r5E8QJkTiaMnb95nmG59RQk2Brnak
P7J8hG8+5j5I/VmYtXCDscxG7jARVkIYnfpJsNaOTaB/yf+CBADD7yrwpPqigrGE
abPkoyuRJ0OypNYEF65cxpq//ZcukHeeDJzpE6vdoW71eevN5CmqHcTZ+LKti+vL
IgyjAuWJsQwsdVnpCx8MSF3DWl0Eopd4G5Si14S35MxztkdfQNV1q7RvuKaeGpnv
vjJEo48m5HNhOtwJjqbSWF3MlnubwhJ32kvYe3mgXnjt30re++396/dA694jv4MV
apY9mI/pzk3uyhnCCxAu/UGpzfPIVgE6e9P4UUWNk39MprW4mkJXSdPi4afw8OVu
iUI+gTW6RLsIoIOoxmt1DJl8A13iXRohQaL7RqMIlWBe3gzSLkco1/8LcsX0xMxP
Tmq1O0xauyi1vxlcLI2J9QyvmBZLMs2EKOgYUdv7QGgQD1kdBWvxJeK44AzXuTuU
4aPJCr21qF128MsKKyOYqfDPJFOZqDg9mNV2QNgDj1mcfWfSgvLv5krQJyhhGlgL
Vhp0yzPO5pPDFlgEMn/ZV+8PwEuaKAanYzU4fS+UY3eOGyZqgTjDWBtFZONKKGvj
fAzXi0ebyL9W0BovrJhIYGOs7akaZKopARnuzLrY7hU4rRRaa3IOTrtgyM+wuwvj
gt5o9l39RwKxgwsu+vGwDTXwxr6RLSqnvtnL1YGgngbiGYiEnqcgzeQib/71sXwL
hTfr4hiHzlpGqKhxLJ9Z5PHKyg9WaVx6xVVVOK92v1YYT7/4ONbEY66a99ZO7r0u
eXviKtkFZghlMHqA9EmUwvbkQOtp1Ta4+QI448FQn/pZSKIom30wU/OOGqp1PETG
H+3PZvBcN6V3i4lHjUqez73MaYLdnt1QYYELH1SfiG7Now5vzOamEfVyhfi/E4dH
ncAb6WLi+zFFruYBMX50hRd+b3NJH/hs7IxbqCF4gDlpphHRTJgtGZvWpykY8MYR
/7EBIAf+kV7XdoKi+xzW29axKhuE4Xs8L1jFGUYhcYh2BEL7dNijeFdiugHg5lu3
Ewyb6+5b4ZZ2m6DF1L3GIe/AMB1UaD0LWOPtQbEjo6Sii/2HD97XEA6nSTONBMPO
XdLVVJ9Cwch9v2N1mojAiyIcbzQx5ewbNS01OJyzbYq3QzBy6GayxL9pEQ1sj5v9
4vA//rKPX8+OdrK2+UzQCSOHgvzj8yVTPxm6h9fyX8ns+LGRhe6FqEyp8gafDqhD
vT5Tla5mJKlgJjgIbZPoRNJjIoaISyHx2LJYWHVFOw4NgeVDxwMhRUBIU3pN8UpR
BQQDt98yPdngr+3oO6GPSYrgV3rMvlPJ329rssc4Sm4kBTKm003ipFNwvaCcb5q9
9JemzlzEoX1q9TeaudBeH61beLWPTvv3zQi+ep2WmXgfwCD0qFkQRrTYNv6d81lf
hDEi0DoxNfHjZAjo81UQ/5Fpw+UaqMZsPshFhs4e1aU0MKnEfsdiebrj7x2Ny7Kg
Jb/hubpx/LeKNet03ICqsLwb8/TK75cLQHWpDfdcYmH+AhDqzhcd2Z3gU3Xfdwbc
ilWI37FRJFRplvGlXxmwOfvaprLev4q3uJz/nqB33Jtqjwywi8IlhZm7745SzUmN
68ZzhEmaTsiaOcFwF8f7Bo+rTBrx29dEtg4lg29xcF121hO/RMJoB1Vi6xitxJHz
7afhc8fe6xHHrfVr6eoB8AfQA22dlZIFpSWpYp0I4wxm9W8pO+GmvtvTL7ry1XRB
TQgL+AASQ+7ATA/xl80uNwlMYx9eVRQbxR2+pdsOpu1xWT+x2tGWo4cKSg8SVDLw
U1s9MzJsP42ZJVUCC0I7pVv8IoXmUA2jj9Lz9BQsu5JPWMdJtIi0WgqBkvzsrjLt
4ZX+WWmC+DmDtmy1jv66BukeAl6075ac04Xm6eboctuVSHrV5wvW1qFY/7XWcfu1
zOhPTQnxKUgS0HJmDc0Q7w3Bp6awraQH9yKSn0k7+WqncdS7c9yvJK8OtUZwMPfr
yAMmhZF4f13vEOWcZzqIj4qbhiCmODnauknQFN7u+5ya0yiJBgLiWTPbCNq57mH9
XE2CgbLAS8cNg2CGHNVvU4dPxnNYwXmjflgEJUS8D0CALaSFaE+AmacPQwTZrEeK
sEYo+Wge9gWNFOS6cSpE5fXWOMChQj/zJ/I+ESm6McxYtckmY0t6UWubVnQ5R1Go
gxiL/wCTmG0ofAMG75oTBVdC2GNbd7OfPpFXMGHlnLM1l/tiow8C0VdTG9r+4XvR
ncVvq+sV34Tyhxb8K9OYLSAfwyvstkq0KGPkustulPC7cjtFkNvK/qSM1IdkjUzi
yJuBGruQw+Sz65fagdxAim+FbRDDCDgsFblPL1n2vNFzmRlkDdryMWbWxMEb8/SF
qICK6pObKD3yuVWQZUJjpccq/+L7wpsufolV1FwjHfzf4HdxK7H/GcE8IhRB+VNw
BVLcROflza+UvnLY13XGVBWrJplioK3B9BOkhLKQSgDV0uRy2btSzUsYaqD80nWJ
OtP5lhx25FDaocmETXVYyKu1astnk3WntdKWRGYwAMWxkhm1TK+n0b8E00GDamYp
wdEE0FDBqXvgsQkd820kb8Zpkv8XIHZ3l/g9tY9ioQlE/SJlt7ff+LvaDW/MSQsi
K9s5VawIVFjljCyUGEFf8DaELWon00KW9q08484RjKn3y/x963VKEkUiXBqNI4Fu
B3j+XXx7yuoEC9Eovthcf1YCVqd2rreD/Rhirr2BL3gN6qyxHhYaXOFh9Rs9hqLf
C4V8FfB60h7wZZDX9Hin5x8CcfKFbo0KAESnANxhyC0mGWtaAq2uMPgfoSG3m4TU
VQ3tUU8a32rx7HuPuURkoTnHTeqZJYhOv/Ecgy6aa0lrPCxHjtonV9DOwz4tgSRF
M61UAqR+XL41H+prDUKoJ1SCdALcIYd87G7ZaeEi8xO2h3grr451ftOGAdsWM3gU
SrEVlKwOJHHwRC5/kLGvcZGnvA3bnVA1SNAbGbGBZT3o4eVTRfk3BEjtNkGqGtW3
jc4+mYRKeM+EL+ivrfrpq3UpeStmS6kOG5u3g+pZzYPZqNBRWXdtSN+pulDF9ykx
pOqgLKRpFem5RPXihe06nDEi+gr2gSIYj1g35JGF1UxmPf48Vk6oD0gwP4zpcQ1g
g23jEizqsOhW9Lt15hwHNlfcnir5tvSUBsf2eiE1zeoXZxBjC72c8lBKSsJpHHcN
+LG0/tRNGaRk1alUGzuHfhd2NH+O1i/aV95nJFdNXbESezsF3m+RfS6bzoskUJGy
64a/C9GR16l4PQCttkU16cFL4U+r0VB/9z1aWAri3nTwfacaxLpWwnrKALDExBHW
wcze82UA0sypkjXHeI28sGp5c9jv31BG7hjSoSLCuZzyuz6/GUI2NWL5CSvXGKXX
4dKvu9hhLN4NgiACNu9apbrmNhAw25hugiYjk04liF+68XZvCvVP+fjlmHFSCGw8
NYFzcbbziE1tAfD9+OGr1RDLyCPHGQ7cpevzDJcP+rV3ATzN3FetOOjY+yyYrYWj
wY8jremev94VAssWp/N4gMAx2bERvfIQy8YEjL+wAOC9Q8sCkZn8MpuKa2qixm3T
9a/pCrwe4iiB5tx1PgDemruDjp2H1aSJYRzcxm+GrImq1PcBMJd878Xg/GITUziB
jyr+PkyhevOgJuJfHLm4OpOXQu7FolLSusBWxCVMYZmV0dVwWMbMgsDef395tCJD
p2NWTbuaYuWeXGNOQnmV7O6qIoIw4blqzUvFQ474ngSxugDQ7lmG4fII3e2NNhMd
/g7P9ozxojCYmv1LnFFmWU4ywQ2VyeGve4g67yF1KGltVNozSieWQ7RI0QnPAQOn
5uw2F35CN3e/Uyy0YbFxvbj9NJ3cTOPjJLJ9AT19fqGe8dtbvs0COCge769WS3sk
wYt9KOe481WN0ea0SRe4FrxLQmaERnWRbM9GAS+JzUsYAz/hAputZ0BKTHSR2iJ5
Q9EHL5Tv1rHicUDzQA3OEeGF5eJTqhhnBOFPi3V+w3ZnE0oYUccYBkJbblbu4ldF
hTF/MKMrclDI/mbRrbzqxruaBi/4yf2tdZ+v/Bto3VWF17WnM7Bx+DYLtz1oh9Ex
8ACeHB2eoeCWAkskPki+GWPBYM1O+umEhQNlVcq7C/9jc7bdVXRsLaNtexoxuO9j
/T0rcPGimxfR9iabLGRPLr4MqMy+oJmiqc6SrWJxCXtkFc1w93rkcYkNP/SVs9cd
VEWv+EcXfVpi/y8eegSNGHqH97NoKUaN5yctCiksqjtMNFxAXa5OfzihMV5zvXCM
KgCJHlMi69H+DQr15qQ0myllqx4JFkvPF6a/yibWCgTIdyZydbQF02sdaeXak8J6
Pzb/GkM2QONvWnT+dHVIPsCHx1p9s41WHe0aCyQCwAr/QQBET2oiOFupwccNw0CG
H/ujBvITtE5L46FY81JVP78GJy3BMF6ndbb0NlrDGAOqcm6f2qaxv9cVIE/Lm+0P
4lG2epOeUds1mVQPatBHZVFL7C6m9laoRwzMgFthP9RJRkedt56r5TevxGcMFrou
xH9xrGbR2TnEL6BfvMtvba0M7R7otVpfJkHEws+L1u9Q9VYomzGPeJSHzRJxphdf
Q8LbgxIIFZyhUW/dtLee+CesM15ajlx4GS19xxP/8ByUX2IZPJuOmei9sfZS9fCU
nIwa17tu9NXtV2rhsWQx4+GOnQaQlIKyHAG6UQ+nJHuvfT9iWjG/IQQtAWUehiKH
7RGWWqFTwv+cXeAKkTW2caSHkZmHVmYmeJTj4k5Fp6VORaO91O5lAZW683DZTIs8
8cqf/QwM1eiHu5YHjvNTilLth3jA5aFghBaC/zHR60Lz3sWH0hX9etCJs9oZrFaJ
dFAwGrclrSGEqNE8LYmeIbdPEvzjQDlTrIRRYLOHdj13pjqsOwOHUHz+J+SiNr5B
NuYm03g6E2dji/AK9jnAioZve4sPE3pxPWW1IjwzcIszR2AOPCtKcu1znP3xXPiK
Pbl3xN+GmsCH08HeUqPcB9beLP9isT6aFu/cq9mzkqPRxUhP7HC3ZN/XWyqOHMJ5
oReJe2Zcnq6LADM7Vau/JqNndHLThggs19DxMDzv0ht8Xz1XZI9ZPhcHj8O1wTGH
oNN1Bfo5fwb2uzVYzerpF+VJCe/WoBghgMNYddihCnID3CxmOpKRa8vjxUyewPw9
MCPyr4KLXopZOk4dvTAfL/P2NBYfNA9/ixZjVjHAMbpKLSEDEWesFNX2SVF3MjsQ
Vos4ZRYDnV+zGAOIHHi1nUjY1wL1mJMRII0DNMScPRmSsQH1WJb7O+ItnvoggYP8
9cu+A+7JupZ7cfJCK0mx7Lwxgzna/AKtg0Csq91GDShZVuoX1hh3Fzl3tTUouIsr
SVOPUNVc4NmeGAdrbE1mMEtBgAt/B4KClnjYjbsl10INXilOP91Kmp23NpnPpn5i
euaMxBQl7Q2DIL1PJbYxqGnKWVnZcp4raJcajxW1yT2FY3hCToygt0P6UAaSMtkP
iRmf8IOHzE4bcXVoNtmLerumJjNY3G11C/Ur9XB08e6+AeT20HYIO9LVSAdjl+Z4
FY5R9pWaqj1XG6T992Ir9Oe1mD7vkEWBm01Q2z9a24Y2QWS6sZ0aLiGyqVeFokC+
Ti7e664q8Acl01lMuLIFgjMWDpS2LR2GLiSUaHOZtZOhV6pPadJ9K9+uUEJKr4rN
e8Yna8eOQTaEljk2N4LHbFjj9Xmuc8qRLHZQCxud3YSmt6CCQfavWod+DTunhX4x
/5oR3BSnR3gAVYHj0ggANw4qPDQvYmxfxFTzxuh6Qs/blB7aFXk1R1r2VLeKZ+N2
vA2OmSv95BTLVNIabZqheKaxleXZIeiirv0eUaSJS1GdFR9lGnX0/XiF6WHr9mAt
piccpJMnuhwNSNb2FoLhS9e4+QuSinVMcAvskMpQYPmj67ObwhKWy0gdcZpkan42
mxWISfREFHeXOmFn7y57AGwgbt984WrGTIYIoTOjlwaVheCpy8ayGiv737KuA5zw
+iRWQgVGjLAI6KwGrLKw2bg8zFEBRQOICveJQRLI0puqlJOW8/J6/+9Rc1AxfCEI
GnfbIE1EMfNZsfFgUmnRJwf8IDGX+MGR7RX0STqaFCQBBP8Ne2saY4q6msGkAeMY
k2vPvdQBa8qM3Hgce6X4FmbrJZ7kjqHLmWzmitaZiRO0eTAPWMQqTyk4Ym6Y19Pf
Sn9ULDupPSy6hB1UxOM4QHDOeUIZEiCGBJPvBozaXVIa1q5l2AzuJ4QYQfemuoxf
zkwyqtmEd4WmwCsaoV3y3td7uUzO/e00X3KfXNn8dqXAFmirNtefpdaPORbHyE3z
YafXaN8dOpQIvlLjnT6rCHaD0mnhJuyItO6IRQu+C77KjeObaSE3PWhJrsFKnIYj
fpLm1+pzo/Ke331P4pbc3vjsopzt8vBuYpiliMpk6FX4f9nQVnI0ImozQhJDXO3P
eiWdkj5Htvf6R5QDgCll3Y2mGXgXmxAWB0MeV9EwewnGwkYTzo5OqceRGyZlJAC1
uYN1PQeYRPKfjMx1gyGcG6bsapSAjgvIhc60xW4UwQqlgJlHUXCash3MBeEUZmZY
4PXRTkTIxSV0PLxJ4x0fJ9pj4Kp/pmqX+qcOVTRnP8DJ7qp0Zz+ya6AEnxLG1oJA
xX6JgLcvLOEJxtCC2v+v1ha0V0fX74P0rrUDKthGy1o2/7FegnOOiRp3oFOJPZ9r
VJiYwZNfaQ5Hx4XS+tzuH5sU1RG3Fcw5OBN+mrFbsMlxbnjycPnVYQqgefXkZftd
JTLV8XJTNjawOqp58u3Vmk/q77eHp3PLdpxWHcLa4aH8phR6K7qb42bClThFIHGB
tOZimtNKsyWQMRfatqCSeswWf4ePbMzxyEIZACt29T6uhHZwPGHRtyc+JaplQUuZ
a2qcs+ENncyUQxZWSRAQFsAzqQtg4XOMDMtLRh2MGGm5drdx5geQcGb5shQUxA5Z
HYccTmC1tuCnWk2GhwXrjcjKNlgx3nwiblrSOVi45HRGbHG7LE1wTqtGCfY434jt
s2OtLw9EugGcCEPsys6goQbwRHChinwLiYF4fPy/54ipGPHeKXTUd4l/qemTCilH
hWiivbaIdbb/AjA5f2OqrQ2Ictd5vu7Xfqk7N7TDxg8t2zTUQ+j6CXZX90hsmuno
edp0w4SlZsQ8M1gZbjYNcK+jq9qNWPlgqiUnBxNmrF/poyKoH2Dhyrp/C/MyqNQv
fbvkN8DrwTnZQ0A8wcDPvhVVve9CCE8+Jvp4/9m9EAoFS3LvkEa0Aq8AxOk1RNsl
PKPYtMiO/X1BVZH63iJjHxyMaAcTR/pppCJ+Nl9lSqeYSrhONXIbT4PWHI+g+tN8
b5BBJq7/HRN5T+ugB2/YztDQYS5WPq8bmmX09sZuBDYkAM23qcASOo/Y7Nbz6dRA
KwTK1Dtjuqbw3cDgIuvaGBjkl1H4uzF3s8mQmKo92jDIexcYR9rsWoGjkaLVJzdm
8ks9WozsIYRlqf+k5pL8QYX3Tqj4nILaG39QjH5bBGZKkukaFgHgsIgtmXeMuzfR
78bij2jCEb9CqisIjzDnsp1VL2GtpT3l/bgZrzN0i1rX0MZO0md2jRMirNc3bpT8
bpf26rE6sw9l2Gc24SkaH4egK5OwxBBi50hB0lOwZ/liXRYjeagIlBolyA5mnnhy
lgrYgsVCoHsrECsppJbTRgzhTQeRk+lO4zcwcE7EYdCFZKJUqWtuHyDmyHbDjqGV
96z0JhmxkfGRK5ooOIzXxX9NWETqFRRJz/LAyeuAptvQmg2tUymPNDBMI+Ze/aut
GTk4+X/QBF2w8FY57StbjJVkNWJ2gSG3pVtHjXwK6qhdTHOEXnWynhAlWm2D4EGd
W6HS5mgGiA242YHpTMpRFuSXz8ImeWbmQRZ7RLEZmtjrUqX7E8CtztTYk5IwciUh
rZBpMydV7bHsTJs3OmNONgtyvK7PkVsVXPQa3QDkwQxdMV2taruolrubuZiepx3w
f09C3UESvfPkrdUFTnxs7F8D1GrmvkoIy/dUGioc4gqM4uGXLrZKDVB159DVGHoz
rD9R1n4xf7tHaQKByLKwRF6MPRuHZSW5KIdDAZt3yiu6n0JIEUbPKAz1f1I9+s2S
Ej5Z8HfhfU6yS9Uy9vU2qdlA+3NEZeQUE8cRRZCAaZ/4M3y68xkWpbasy/yGG8rx
LvwKpK7wpYKVZQ9e2BeDHm5lT/Dc+sZiZ2VRBVDjEzWDjg/LKcx4szIiKKW3b8Sy
0+fY8aZa1KLMCBjQYrEdD1afa/MJuECMSxf7kXnnZZcCvAb/PmGFUF7IZrH+j4ZT
iLc6B0bqOn0iOfTSmV5DR5mNdP1BTBHb3b13oKlqbc50uAm/4yJSd7WJDDHUEYxY
/s51rg8T1+x/A8wlbfKVmKU/r+HKUpri7w1kKbfHCWMLjlYlWXFuQCSepCQi3gQI
FJt8nWG7pgupn7ouUCvTulhHc7xdUnDrrHJvMA4RYmzC3Qd657cVwfUJJwbI/k2g
1J2rN/O6xEz4KFL2k5w8JBk7ruie9GuLnJP4wbkpO5sQO9yToxBumHSI2Wr1NYac
pWjwsbDOd4cyhsJ1MRIaxMo888jbbT/Ast7KT415Cxv2LVDU6eACWibW1KNfe9Ce
88dkONyZFp8iFLpe3XNfKUQnDPS9yd3K5VL1a28W7zca1a5zyH0k1nCQ5d76avSE
GqBtpW5Pjl4innEEusOuCf7r80UFs9JHm9+3hfkLF6xLsEo90aRLj6SuSEeAtII8
UhmwIPoprDT7bxU13yGpXjVDR6pSjhOB2Kwpb3AeJy3d8l+g+CLcDPN+PhyHYErb
ePUNcQbY974LRXhafh8mKgDCIee+RLap30E0sAg5zbpXyq0vz8lmui8mnG0W7hYH
7QC1X8bqEQ65ULctwCJyMcJJDhXYY8nuGp3tkOh7mHVTPjOjm4v3lM7+qHJAoX0w
nhvqCy6TG6jAxqyfb/rfoKC4NThjUut9XRkPwiZSSLVEtuqwbu2LjMuCjuWQj5sm
flxGmHPMYeBD1lT4RrF9jHWczToNEq9FX+jV6j7mp0q8Nu9Rw3kk44veXaerVRex
ZfCkOtsf19bjvqcfL3ICLi8yDBO6NZ3zWPjtXYdvFy+7jCENHRd6KPfiLJdOA2A4
kWlVdYhGKhmgKIBXLSuNnGcpde0NJ8B7Btw6ipqE3Rccrb/3LBdcxXESPwg6JjqW
rEPyiHCwCsD19WQ6SV0V9HxLRUsf8OZClQNTu13lEvHsYEFcBeAaZHruuzaulCGB
PLDOln9JgZawSzJItP0RsebanLqCmnEHOnyrCesl2ECldK6hM7PkcvCM2nGEYq58
kVrBsPTbNa5Cmef1MMLdREgzArQ1FEAuHJOQXpExIrQDrxivexzWIPIPWqbQtigz
DmfrsE/eoObV15SBeYYtZVuzMjRzsh3q9IACrRKaHXxKDenxW+tQUPFQOEzquGnV
QzBsmHlfXGVXCoqS9X2UhkgdsyvY0wbNxXV+aOrfLvj2WnykJWCAuGGBTyVFBjKi
OIZlVsC/BGsl8Tm41cTS/5eWrQzlotNN7yZs/YKFcLr9x1x8iKDPrW+1shzupddy
YfbI9YA5pKpEFAd70exWtHy/Jk2yrWrqeKlFZfS+FQXbN04TQ5jh409Jnn4Ob/hM
uWlUr5LG9/m0fn7nEJu2Km/OlRv7DsoVsLBSlnnuqaRqUmOV627wlyj2/nFSa+Dx
kNCoQn0Z4QXOhr0nJtOQg9Jr48vu+JZ1FKvR6MzN/BURMdw0nnwn082N2Go4Efey
nZIswS8IsNXehZ/gQJHEq8NNE7xDOy1O+/FNTm7aYfu4A8RPUhHfC9vaJxHGUKQW
mKneHim/kro+KhUJOt49rYf+6j0o0NGzQcQYmBwJIk+p7FpFWTJ5qXPx0ahj92NZ
BLtNhLioRuJOAjiilEFrEBGeYsQ4zSBTlo9spq/ucYle27Qqh/mlnalrskdEZViB
GnWq68ULj6WF1DeRh7KUmr/vvE0Xag8UtIwAflCHxvuI+cCK2vhpgW5ql+7MF8Zv
xPhoqiZyeiGTQTBVsL2+ERIDFZK52TEnst8alxa7dnIfEG/WrnYh3+tJdoOQQaUU
q7SGr/nUGhxydNlaE41jS9jHEB1n0jqr95xsMwKtqf3A+DajcI55eRoJ0cLCWvZP
1ZFpiyTqqHwCJHylHqButWPgXUIxGnHkBIyJ45viyHDy2EKawnYizn0VbhXUfr4N
J8PKeFmH5hyLXhuqBZDgSjeMBCoABHYvILiCR0gBsVC5ymDyrxIftgYv36afraIi
5rGRnf+ZHgKKQ8pK1Fic/efFUpaimzZQvShJhDC/570GQG7iY87KAQ5+NO8ZcoYR
04Q2Pvp0MS/iUJJ6uXiJZ7DDzcHq5OGdd+C8A5wo5USS+5BG4eAiIdf1G4D3gket
YxBS/LCL8MtOrFgc/YFQNrg7avoZxpRTIXdiZXR1hmU6cRyc2DBk92aJIhk8zQLl
79PanBCk9Ep6YbQdC86X53l0/RxtF0UVSb8MEAjcYWGtKn6C4ooSosFixfuPuWs4
W1FZMdZPJoKim30rgew6I3dMUpwqgm1e04ecNweJ7T605PrxtZ+HQTZOkhKT6C2+
aAKLKP07u5fE1PfRh2N4p5f3P9rWDnubSxjCQfS8AvZnlPwASGQyUU2HfdZeJ1kl
UR2k3X5xboe1FFlStrpiK6pI7XrKWYAxMxjMOd8/bm+v0anqlLYEUPpnr9BOuO9H
qfp4kNmENDhJe3aFFdw9i9wLiFi9ViTu5/uM8Bb8oe70ZHTcQOz0cmB5mDbiXClQ
My7bCi8tiMYopAdlnMzTxoNw436dxqTm9IsV19aSPtSBzYYJ4c7nB/eN7uM7Tsrp
RvwPFHNpSwI1XQtOMs/trmq24Q3eKNlA7s7GfbXY4xRCmKYGdX/QrzNbz61BvPtX
wNHEhu4HbedT+g4jQn5PczkmOsbWCXe6sads1UD+0tgjxr20hCJALxIqGVWWZFKW
0AWje9QYvpNGpk1ycyEK7Lf0A81xZOv1YReVt7rEzQG60MACDsGVNsuI2ygNNUt5
W+WxvxAkiDwpiR9OB6N4DV58UXK6y99HAX8yzev1Nw4LvYkURgzvXmTRKlS9W2D9
z5MCdFl+5N1w9Q2WzDp6DYhcX2BP7PFnMRyTnK8fHUeIfv9p7/pQ1wC/oeo7+xae
WRA+6UXGd8ZypXIS5tGurusyJ9pkfdIPZZUnAoHydMNFYEIE3ktW37l8eUBja1pN
e+oVie3jP4S0h5RYo+Jmelk78s0mb0k1L458x1BWhQc7jgLCB1AwVc1I0RLhOgav
1Ml9QQhvVwEsrsj4pJuU8dRGRSjR73BXYFW/gMCDp4ea8nEUfwChZVpLpP1kla3g
S/BO+MLRNNC8HFlsbieFWl5MwUQmkNq9qsSx+t+zurfi/r86ys4sMxPGptpzxpvY
aAbwZe3QJ1AdwQ2K+1eYXUrD61EJ10fgEiUOEViZ4XUQUbikxMPpUgzU5ccZOTcC
AQPwtMHZuV8AGEI6mojPBiEwoqb5FLLICiF2tX6sf/mHRzAPExnn4VS6il67ixev
gLnbjug67bOgxDCMs6KCuvaJrDxtQTLGr3XZKlSN2lCJs8czuST3n9eYNT82QOHf
pZOyEtvVSz5dzjRJfmaxAGncOkWlcjYr2dZMFEFtq3n9zJZ+HbEBpnMeVxoHnrqV
3gYpyTg0YMkDRwz07NLf6AaXfaiIkTNmh6AN/7S+9be4yiVTK05tl1lgAS2X3PjI
aSIywXuJI+bAI3NYHEcAH/CGuFWhvrnxZZJTdpvtWnvI4DyvJqHc8mVv3jfCD5GA
1Pg4wL7SqkTLrsGZVZ+LiNVs28nFO0M3uOIVzd8KmYVNrLqY3wizFfpE7kJBJtAx
YPPqCh2dVqLfCGnHB3Qfp7JLvPS92ddWnuT7W6FonRPLJQ3MxsBWO1v5RTcMpc0M
Z8S4Cw6fChRUQtF7kTK9CPsODm/bQklcd2gutPGDe2Ep5IiqUI3s3W0L2YzrVOdr
+nDaDkQLSoSx9y3KehT2tF215Azx28CIHEWXtdn8CB996ICXvKx4R+y6Ty3VH3Ug
Qid5AoefP+cPjc2CNJtB1PVvcZh05tUFut1k5BH6G4R9SNsgGb7ZbAqWie9zyZN4
iUM48BQuyO8EforDnv45DiFm1EPs2RAHBiPHSJYXu6S+7pMXC7AwOMHlvV1kUEnW
xRnd/LUnSCSuH6hFQaOhYONxyayKJa80gjxe8AWjezwOgGAE2J08LhgMISx5xYhB
UOYgPM/sxw1rmhKAjt6HBKK3ogoOOAbv2LbILpx+nMCIs5r11kdD1vvm3lJxiIJB
5pnd4jBJ/8YBsBtwL+Q4RyMGmT6cAiwuTyLTb7AzaePSA6UWT2ZIxq7Fn8Vnurso
YajgfaEqQSVzzJIJzgh4nSNcC6bXeT+Wr7YGJnjZo50aZQFw+NW0dF0oi2bxco5A
jtZD52rQdo/yo4DH4PsTSOQBiBoEEi8Wv3JMoYcgYkDn8+C/KcewrxE0BBLLSYq5
TKiriH2NruwQLX5fm97Nt3lk3RcVnhMSCdifAL1TbBtK6Xmz2M+GQpqgaccJ8IW1
d68fkvytbPRjJAEj8fuzpsX67d2ORuydsyx7+DvAuBfzrOoaxyOdJs/xtJGDk//9
slep/VbFtEeTP/ySBmh7Hx2ZDzQafFnpO+g4iJbD5Qn4kSCtqj69fncRXjv4BxbP
et/vBLkDvqubAMqn4PHvKicc9hros3dVIWepNsH6d+P2p0ln83ENtRq7wqRyoKyy
sTjn/LPthcJ08IyVJn9Kih8LVbMMcyqVik+AjnbJuxOd4kWTl4InKV5iRw7C2To1
9548cNhKbT/gcbqHt5FjDFGYU3ZZeNIT9ohyWYXLEIBRO+OMIf0VIkjySbJ+TwTt
FEB2wH5ChT3AQbCoNoiOQsqzrignGiuuSrJBUY94LiBqi9EFDz1sW5Vcx9+Yy2aw
uNEUVlgUKYZJ3biztdvRnN+iU2D4CZMSVgSufMkoUZZZYgUJEZPmimxcqWqjbnhF
J6D7XcvjbILaTsxPQaylbyJOX63MTk+F2M8NsZQD2BJLioSXhc7QJudFBfQ7y+SQ
waLumbgwCbR0WFEUy+/MiAWtkn2Ed8cnPm0ZR+LXLxdCLpET6e43DtFnTumkjtC/
xp5DVezfvkRhmV1xP7O6bqmfkpOgWTVfjktzJtKRjPcaJf/53CgpdyCNcMoZhBwF
Kkoz4QTswCNcsMeTfSvBy+pwrbHVNZY7aAseT7VfByIV7H5hafiDe4RetbmlxOfj
EeIlIUtm3unLD5eUr0YDOe4L838249YFZdl3i6qpbfTkmpkLMp0qLlJVTsaLP2rd
Tj83qqfK6hzVR3iM+3Ux9BaySryFTYIGXvhrZTppfjiMZXc7uj3auRm0Z4ds6Nl2
n/YnH5T5LL8qpHwb0Yeq7yiaJXohI/cBnfDPvZWrtqSyTlU3rQci+SrKNd3ywjvs
BOdyWh7gw0Gz1THXMuRfnRqDQI0lGyYqAevEmZqaHJiU6jS5CGiE3QHaYMdWKTv9
EF8fOoONssci8MJcJAWvJAtPqYMcNklGdSHxu8ENo7ZV1MVsPX15rStktRMAh8Bw
Fk18Hv+zB3G57vjIp2A6J5ndys5jpLDE3yQiDCZ/YE3W44bImWCRxsj7n9YvgGAF
ZJtuabKLFQ4W+vfYamPZq311GmkbDdEgQ93fXyEtT0Povt1I0D86L80+/0IyIAjR
/OqbTmBg/CaiEtHwIZuVvURcM2xAor3PdG4cfKNfLMeaCzmrCc4XJo/7E6W79LLY
a5M+FnRABIu4YuPgqSG+QgyFUTyCcM9Y8OCD0PUQJ+8hElCOfFSh7KT4MvK7EfIK
OurqI3NGXtSkxagtld3QxV8PL2EkbvLCRtuxlAWWLjetHRk8mL2dL9s8FD6vD/qE
hWz7DBgji6HsAkC2sfsPC+WQZFVTwGNsSjPIFBWjoY0o6wNCWTsQD/0W7c5KX08g
LV73MnnY2G9sz1/0XjO9NzSzOT3ytK5F97SPZ3J/95lkDcaEKOtuxa8J/J9uuNrM
s838AKLs6enCSHaZJQnrjY3X0TP+hQozNkQxC9TTldsZHbw7c1U+0q8f0dxYuHJw
qb7286rDWno+D6v8SOwFlEUf2EsUB6i79dSMOz9Pqjs7pmOfUt4wkW8P8yGJHR6S
89+yK7qqTpm2H2MfKDndUJYqNhB2grt2AyKsr33csg/1HIp9+7AJ08EdZt6DaIKg
nbyqyJE6w0SCpq6AMnTb/qYsUmFqH5pUn2cNtac3V+p1NZKu6nFfPsaNwd65jpbv
SnfUjrv/xzObNgmd3CR/fa5oFYHPJEwQC0l8cwOR1xtWpidJzmt0StUrDt5dF7AA
yK3A5AeJshYtlTS4JB/fQsO6KHJbI8G5X1NwUZv8kzHabsXXo0ugbxomrivDu9V3
Gdk4J/o/96W4A4e9BiF3xEN8GSOlth3SFvBNb6TaoPaiwk9hIBIYx4bmBPQGCCVw
uYOkCcdLdP/X9lSmwYtJZxKc+DvNwACFTSV7qEJBuxNVIgyLT0lXY1D1/clDMbCB
8cSkhIL0s3F8q3gV5noDIzuB7/0Ee5/qCfhKFBw3ep25BeNOJbo+2TxYN+efb39+
C3xsTIZq69YbZbG5/HpJUk81tsHNPVEKJzWcJ0bRap6d/k0z0f5Lf1vqfMYgiF4Z
GzsKij7iOAMvsleDbOmyiSE++si2Gdhv6de1PWqCZaWvgh14z3pbZYnMxsH9lpKu
+ErwSp9msWZBwicTHsxMo8OQrdGgEolan23vkgMjBzOFXH3FkQJb37JWyvVnwT1y
TqFLuuqh604s/e/gqiCFtayWnfnGMBwGqaQRUWqCbn/FxPzTRwPwLol5G5B+AVU6
h7hjo2j9uvfVk2NmCflzsdH4BfoIk/62RiB1Ld0BFT3cxEHtpZhkGb6vgmH8rgbL
/fKDoKVcbU1p/keYKIJfp/RlVxwwk8/uC/fugGVWYcTgYNPeCUaLabk73/HDF64V
Ube+wfrypJHmWtr5KoHGXb8zGeufJ7byplQLNly3kJHn03btSJEiWeSMEC/3/1qZ
SvHcfkdz74zZgRfXq6F2wkhJPAIt4CSX0+uD2mueyNmYq4heaChDLGXULcbZsRhP
zpA87AalJn2m2dtf4XyjhnPJcnwBBP13ogMKfxIImJrrlldtYaDqaC5upBjgy0g+
p29IRQOVuxgM7bb+l9ZH5m5pjVs+9Qcp4moVbTIv8OLk8mga31xTTpglelitkhRQ
gVRHsryz2Aqu6iYmdznrULh5ny3kv+ks1fQ08vHVx9G6WEE5bAjdvWT/KUo0rrdc
30LJ/DGL1rugZqZ5Bfg4BGFQX1wCEfX7F/VLsKlJmxYUqUxoNP1xuLOzc5wo1kOA
DX+4pzBdp5DAU5LK3epJv9U4HKDbLO40X7g2ENhNPNcZQvf53aSLHqPOmL7U/hge
LC3jMZb6u1joAZwKT3y37wZF4QhQatpYRQxTlbjWHTc31vMVP4VQAp6ieZhWxe/B
CLcVYVgKlRuuDq6O/VNTR+kRaUug351s192vjCOqT5G64sCfMgCIAeuhmwVM+yPe
b73Ow98bfAJqxi4t60XTCRM29X90ZUODeQFrgS5u1YhGCapaYp1cksyFc7T8tRBg
7Mvo4pWXiErD7DtNLlxV1X11kYqTa9NcLXIRtb2/uM74WGNi8Z39Yhp1w8mHnUxb
pIrX+P8fEr6WEu13y5JdWve5h0rGWEPbiVbhv1j3Vry/68dI4Mnho5OxY4/+a/cq
MoncAHrQm30FXWzGBJsYZaZ+xt4OE32P40Htzc/lrNK+57sxt/wjB6I7SwEPxmHQ
RnDGmdviflpxkMXarYXoBVNyD9/lOJ2h6fulr/PEKho4vWxYG1mIEsZzPgjhyJJN
t1x05lUwz2g+7n1Z/c9Wxecx9GdQdvnjPaW2OpY1Tvh1q0Syx9zZ9o3alC+uQM9a
tb+rAnH6aFSipoBwA2ARmDLFDjqZodzWK55i1vvQlS/Sg1SgXYeOiRAVl6lfs2I2
Gakpwl/Tr/Lu9fgOgGwD1H4YaWMvQ1R7HuXobGV3sTdVRc1ItJLde3dW1QRSIV7m
0sAxxSCFYpCGMHazz49nKKwIOPPPZ5OjQpO/GO60Ju04/zH6Hp5jJTHd7zfw7vP+
wNpoS84kevG1j8kUOBdeQY9fklXoK1fPQ3lzgnmxkNm7mFbCTwetTS1cJRUyYr45
0wdp6ACmOEWKLzTeTYc8wyUexgUMQBS8Gn84gS6tEDfxEIM6guF9PkUCCpIQl6ad
57X1tPEFErNc1IZq2U3zZTjy/rIPAopxiqJzVdAxfRDDQ+8B6Pu7WQ0aueCE0YzR
FiLdjw3uxfztXh6iptT4i6VH9WLHtjnZU4pS0nprWpqFvx0JKMT9JOjzCml/Q0jG
47LJzpQeHynqQvFdZn5Y8Ajvft43OM1Xe7neRcjZexvz9LZ2gMfJmeL3KTTIqb+O
d2XmmuMFPl1C0TmKm21lhlBnUGk2NKgWc8lg1DcfEA/AK04tPmbvjZhYPqcA612F
tINdLBD6BaLB6AdwGKqNi3PSenrX2b51wxRoklOVuQyzzxzyTOKQTw+vzuHouWvi
jbWdQx4dvyu5l8pvoJKVWSAqXQNY7uoRbv6YD87zIgfWpCleZqqIIb5e+MpEiEKR
N05zVRcTDIe+uzGiS+LPkg9d5Lq0jznpi0zDE3+1drjm1zzpMAOlsBsdI7ZJAvL/
n3lDLoLqfca/GRCLqKWUJHQr9gsGxOVggDShjgiOBcttVwgLU4balJrxDhQj1rfh
4st7tY1wKT5LKXbAeVV1uazRGjzr2ozSjRzBf4xgZdx2KRLtnDFhztQzGF17iBBg
hqXRQKYjnDwoEFV+iFqqcS7GNK+oNnT4I+xc6w9DRVuMWn+xZH+d9LVMIY9wQP0Q
A1CKM/iXoP0ws6pggnVhiWQ7KgCOeg81wgRbdlM5RqLz8XFNo5KWiEJC+8Wua/xL
sEUdLP5kSBvbAT/JczZlwMorlFOIFVlGOSUVUeIkaAujvE81rYh9B0T/Sp6BDSM9
OIYSD6zStT+KKfYDwFeE3oQuVRmXZcvIcd5s1BhPGD+RnUZRx3ophGk8txQw8vew
iav0rUXvbntq9EkRFMDBGaUNG502FHbKlnysBQLbVbjmPrJcHIK31mW/bOq2Tu0s
lb/B+hee4E7EplSeH8uNGZBoL5Uu4cFwtYnu2+cqVUqgFcsN1ZOvRicwQztkIRY1
TUywOoo5wHagzudcWpgUHvLRb5REAC3uQX4ZLsZ6DtKKg4EoH32cPbdglU2nP3Ah
plHn8lnW/FB9eKh5lxD1Mq2ooIAQG7hfqkj7CLHsHjZGSXIk9cMKJdz44U19mBFW
o7av7bPQosS7/nhye3o6oBk9L17myKRkC1B9VP/y1Hp0DeGdnhupDG+aQeR7M0H7
+8NxAk3ytSishD3OWo907iA3D5+nMFy5DYYhrSfIyJSxw+ccrLBnYsPJ4NXrCILt
EtCRJTjiNPgzCEYyzyXh5esZK5hyOy0CypZ8yn42cyXzpC0VwdS3IbMvY52INMaF
hb3iORX9AdWJXxEAhQkrKISEQ3lrLgFhv1/4nNvmNSBs4RFL7DiGvsr97qGtM/79
ZE0jWwtRoQOn1ia1cg9fKPCRfMg2+jZiaJJctjlIFL9+DtxQMm3n1yvPBl2GfaDk
9sTY68nae44t2hqaOPXPkCItcsJQuDG3D1Kgo0dv+1Jkmu2io5kfcVdRJEPO4S7p
Y+T3fgZcrJ9yKlNqyi4ElPlA9MU1u0AqqrSQok9XmlQNGyS/BFi00xJjzUBNom36
ZoJvlcKGBVbTFbBlnWSM+ozOImLt8ufsGeUpmkodjJxm4ZqL/q9mVZ/M6L2OJYSy
EQXV0v0AowEc2SympmJsifQ8YfED0zEXcG7uYIJR7YIeITybCUogrX3jCkPIVD03
RCG7HG5Q81c5zOjSPfYnXQt/EkTU4Gq5ZaEEJpmnIB1qy0AnTyoxuNEhLiHiQU+k
tiS7+ZU8i7XMt4zXRoZiaT78uzBTED8ez2u/hCWt+QsH7HhOXmsOZJTMwJeI9mfm
5Xu355bEyKIZwAvawA7viJMS5oGoMEcuMj8okbZNseW9IrI9QBd6RQK07Y7UgPYU
8YRIwu4AbKlP2uzOt8ZWVaDaBoR2ZT50MIWzrvBT6pZR1Pgxc07q1odTS2FzZit+
aAQNoJEEqC5cG/1YSnQ0y+4/sn65ud33g+ecF6bMzHOMtNa7SHzCXUBRf5uXH0ht
TdXy/dsxnjvDy5GnorxOcuRZoU56CSp+7OAiwppjUs0Un3C3O6mEiLTyj8HsPiN7
t3aH/9XnGXzAsiK3PbVJDdHMOB1kEQEcJkBIYuQYt8ZrGw8UCLL2GbT4XJoNKb2U
/DnhvmPdY9cGxudZUbReMO8RyWdwb7pXuRDj8/NQgGMV7c66ER7rpTg9vtYHuO20
XGIPsDH1ifMEQHD32hR1jE/LGVmTNvqjzXcnO/kV1FvsRDgy/xbVfhABvDSTLIYw
gark1HiPt8a7De0h+WX5nnmgldIRoafDuV5M0A0ZpZPvHg7KE+dNs8Xbfkzrr0T2
K+wU3ycF7pNQ21dha+TCZX6Pm9rGBu4R7mp1U+53AxvelM7vdCAlcYbWcCzqInZD
ZjbtOqwZ5Cp5sD4ND7MRuz03o+A3fKQRA3qY/0ecU31+OF7YpdOzHRghrhxH6U26
/9yDiQulD9PirLlhHc4CU28487izn8DWSmbuO9wBqKJP1jEz8iqb9Z38ELr18gl9
HX2gTZrt2F3L7TKE222v9g4SuA0RtOuFWZEIz9/Be+Ayvye+tdVdaKP/I0k6jCKi
BtUDZCoEnT3fYP8ullrFwDztUjpBpp8rp1lkq5pSEVnf45ajZ3NWn0hqtC2Bj83M
7+BdkQFzTu3huNMexkTr6dsbCKsxzvIL7aK/O2G4IPHQgMOnCV0FxjBa56y6bpv3
2bQx7QqZL42Zz4GTPBuG45y/HpQVKjfloLDYa3sj3Xbex8zUB++91tDZcMOSgfIe
2Sr0VYvxYB+3SbsuPqOEYR0CUkItOopnXTlgcClp4453My0UZiyc10Y4J5e7jJCb
KjtUEwrq/P2V0gWVck+c/hRsB1d5F5Gz+rF44b5b1NgsPoOLzXV8hZJVg1r3/oxF
KOUmbpxrsM450s4iMjSRD0y/1r2eUqhrXEibn7+FfALwX15/LPGl7ylzGbfntRHq
HuWR3GTPGUylq3ScooMFx/fIm6bHg1PvJtwolmMrrfSngvhcFGFsA5mLNebW874z
NibXca1sds0RrqSkoC1+vMnzfE3DkfSwKSax/Ezt2Y1P3l8EYt2jGFyzxKZgJBQd
13GF/Xw1eu/bfLHQ6tNDSz+RGvfCE2/r0Qub5B2ZksEFC1nr5ZF5bGDdyon0rCCf
m7/ihi+695PRLUhNfkD7BkXAAJ+J5zFMS+u6l7f2eX37rWVelx9fbYrZ1Kj6Zkcd
jxNDkd7NuIPZuK9IouVJW1XgqGIMEDvdj2cSQLRXNJQw8Y47R4rLtOY7uoWYCyvB
d7sBDdSTR4IYB7XlKZD1iffrlnenVmIitEgodVBGM2MMVKzLTvn2WU4IYf8ju/p7
e1OEPHLZE81RNp9bbpKXJHgniy+TM7/kEcqeP+9F3uaxvP51OECFkAxa63m04gW7
uH4Tt/cOfI8XHtgG1NZJzLTqP8ILy3KsQStGTgexGxdKkSFaiJRiZmg42YykjIqF
fQvZ08S1S/GnbOOjf+woKcwZwCYeENmMKVvt6g522r+/bJPUnd/V13CqkiAYG7Zc
m6lT/vS/VffE6GehdSB5Qzzk+QvlkNH+JaRKYnQ8MaYf5mt3Zozh31jgc6L7dYLP
DIaUwZqKRXA1BrMkaGfkTvPrqsf2065pvHVsc4e6FbW3WdWwOYMs3YKccvFs+w8s
BQcerjqacDWfKOYEXdPHoTDeAGD6Af8MOxqOSiXaggEj2L2dDGNohAFgtecRItlN
LrXX35z38ZmZqVyVsStdlnxyRH21J9p1njUk88JyvyQ796eBTOFhD71HKZasFLK1
Vbqpf9iVAcaTfyOCUX4OLknSiA3LZgEEhqaOth4oQqXEzZ5zEJWel4cGMzkO7Ucl
X8j7lPLo3S0+FaOnsAHrHr0utNwCVleZN5RLm+55YXR3xK+mUid9xdPG0eYwJO2g
t8yPsrWG2KIumV7/ljZF0aOmjYwW3I9lJ1R+mpB6Eiql2i8RWyjBN3gGWKu3PiFH
D9r8ybMTd8VA6Z+Vpx/rWdZ08wjnu3rHnk1bymPo1agi2SkP3TMttL5o0WkllUeH
j8F+o/CwYbZktkPQlDLCW2pn8TFcZiNzGI9p+ishLJkJnBpP1IiD1r7jxt5NWza5
oobyREhVELPuxcjntbcoMaR6bFpN6PRHoKw+rWdoj3smBN9WssG5Qcluk9+SFhf7
Kf4Q9BHjmsr7GBTcBn/D6H9kNrp/qAptyj0vmUARkYontmNLJwgunTjSqdycTKjK
X5HaGXXXJsVhdMr4Mz6zVOfLdd5jUN+G4vfrBNWsgNGrhAKSaQi6npOZ98DkI380
Ue517s+1FsdMvIKUQpsqIL/ta1eyEL1kh2dTH1FHvk6rvq4D8wwuzDSrCuHJbvNc
IHR/bn4WPZe60HVXxeBJeGW9ihRY5et7bscx44Sm1kiLU4kqUGAjcGQMKR1PvGwg
seGhlpJaZRzHCNVzhuOboEUP8H6I6sSv5GvwN3YdBqlByKnv4YrSsdyCsv/PPXe2
a9s1NjIuBOrjejbL6HlDNnz14L8soGtch65zB7WgfM88vL8U3OI5jULds1Mqx6tk
qDlrgxBuGIlVib2Gs5VnPd5ghV36xX44VpNsL08NXPkW4Vup7TqdfasS/9vgcmvI
SdQl/4ugCtM2kEu1ZLfyYK9WeNI2E8VuVySOZrloORIKwaIc3PUqGEarmjuEMcHH
aVVq9RCogC9VxkjGYrRmFbFkQpKtDFgBBSvz/0rRuSrU8K+ph4L5JrDoeCRurR1Z
pI7nh2cBHdxEP/RftY+U7Y/Vp8oXzx+35TMnZ9DBmq+YWR3RlzcZTo3kt9yIPN/4
ZM2orYsrWRdXkxgaZhJCzAr4eqwv+fHTPdpAce68xEFoUQJkLPhJATvZqOzjdUpk
nMyyMITVVAdXMLWRAhAHfw59UK7SROflWYyUFPWvL+Xbt2SkzYIK4WXMN1ShDTv/
I8eRkXLD+sfTT6jLCqcVIgVpglPtm5ZmIpEpXRFqPC+vixv6s8GIWO3uY2n13OEE
CANiRZ0fZ7PYKbWmIfb5lt8ABTsG+OngeSknVhC/QDbQf5aHf4ksljmNeToKdyOm
eh2AcMBg5UAEf+v9v95ZlycSB/sO/kC7B9TnHQ2wx0j5cdT6KgME8fQjdYjrykKD
7uJQQm1xecbGa7cP1zipXvs7hzMMC2bgVCeSq3Xi02z82t5nd7NmI2OyjGQ5OX58
yfpy1XFX+SOkPxleJk/MnNBIhnSex//djcyxb7vfzYm9GtLIT5bAAYKANKqEj1Ry
FPc5GhNB1s9wA4QtySosR+dPzlAuBHJLI2zPLCR3SPwK4NxYE/jYOwzdKYX2WoT7
W6SZ4udR6atdTAc8nphcBCkDhqiwXTfUnafCbU93gK4EO/6XrR2RcrpVliSzoOkG
nEuB7mbDKjig8rCC3yewBQ/Xmomat83DZ55v2yGPBe4w3QB6dN7pSj4C1Y23B2pb
VoSsydj4x+tDXRZTsVVarakdeo6hmqic8j6z/6AZNoiKCxxzfUmpBP7e4C8tkSX6
6KFSaSqhxUTFrps211eKQaW5l3LwnenQ78Pbzskz4LsycdEwaVlhB8b4eAzGv4Ff
K1XfWrH0Jo5V52ztsPrToYfEkwdAB/P9E1CxQKNjv3I5fgEcMXA9DNn2brPOX9qN
HJP6o0v87vhw5LRBUEvmfh8/K1+BcFSIU39BdqoOfb2D0uObCvt1d493VW6erXAV
aMoi2TlocDfvouFd0TWMmXkJlVRs5ImCXNFpnSY3b1pOrCMLtWevXSZtDCScwLTR
p5W5eAzEylofX8532MaCdPUS/KW4ZojsIy92/9T63VWbRwIoSR8BtNgLDOBwxXQ8
GzcdrM3rXro3QRXNaORnQbcSfReznV68aAsd3cFIPHEkUT+UySDsvHxcVLBSRhbe
REFeIEq4MVoeH6q2/3Jl43zs0q7ier3aCLsz4ApHkQPoMCoD1/vTCJBZOvax9T4Q
3n7I+jmBNW9SX5nfy89eyhVmFu0n2VN5WeqIs6BL68o1TwmKbCTf+ayrGPpYWhEd
VNlnuUKNa8sZDjvcdum3XDtCLsujXP03Y3nf1nSSYYmmpS6GSui4hrgr3GexNonD
13bIymwI8Aj/wH47A9/+hj02UFMIJ6ugdil9f6yka8RlK3tNA7fBnA+EAeA3AgxI
WhUSiYLHja1a4t4YSUid1nis0/X0UyIrugSD4muIznNY6yaTEoLweR3WBrkYDsE4
+z8rw2Vpb5Cny5fv1GktTQ6km7PxrWcmv6C6ykPpkeOEppUASoUicnNgnEVV7TeF
lBSzEzWgHR1ooCBRbZODTiKdxNdhv1A4TPut3LxotIMxMYQ//MHM4gwMdc4QEdce
kr9DPl9EcxY17wSmbUBlYTRPUs8UXbbGJzO46NNAb2bpZqz5bgSsyxF/A3i13sh2
5VhGYeohI+GLI80Vbq2z6znuNn6lKxco8MzQMpcsniY3dusWVVWb0reHodTA3gDu
btMa8Vs/urUeAmomFt3ZYmO8Gl8Zazo3bdnp/aUzncX0bUt3QNOteHxEQYKJs9cw
BAqZipP+Wems6VADm0PnTUB0maBAJB2RVcgclOHI6nqbDMRd6ftKDiQHDwSQSGAH
tFz2mHIBrG3h9gNKF0QNqNuTJlOrutXEd/mW0mLpAles7mgTrdHiakahsYm63vYa
K8zm8ftYtIh1m+5TANODqb7mLpXqOuQDYLVbalSjW/EK4oDeGI/jmKX5d3MydybP
4/Jgs0hwoRNr+MP3LmezhUmXWhw6bFGjyZxZVMZYmBZtH9yxNk1h8Oc4g/DIpxXI
OX6C+RNUmOGlBZ1C7wrNNpaha8pt+UWL+8tJCwWA76enk/rGcpMsWOuFZgZ4f8a5
G1oQ+UQj26zAmMNFyuJt9Ay7ODr+JXZoyLBwLqtSq2GZPlZM3FbF9hpR35g0/3nI
Im3AWHl4VQHo82WRj1SeaZWICujKGKOiWH95OaXFblchfFSqmQ7cDuDOaz6jNTyT
rRy3FUhXqmWCjUlN2cJMukUPmQayFMZ0M9ataS1B2eVzvc5YbVIj2O7m9tgGjQA+
dS7zwdcIlZI4NtW8Ai0i/S6WPBqrmzcSf3HUH6HJdWqMWPz+XZnYvarkX3Smrp0x
j1N7+DxrFatHSjWS8r9fP9vcsDfLT31m7d5PsFXqvjEolloulibnPLogNJX++xQf
7pSgiXc/etVOWpGHn4xdU0V1lUmA/D4UTiciFfgY/3pAYEHKp+abOis3cF+qP9qb
7OvF1MLCqtlHRP8D8ap9z5GpIm0FNJf1ihSr6KIoMpLOi+7m8lPu8nPGHChukAS3
kB4sAemJYOW+NBt51lE/vnVsxz8cq1O11yEk6hi5EsArKFVtIQjRuPWZsH37C9Xm
g1+cCjxRYhHaVf7KV6fj4Ax33LCHf3Lh9mITPMAvmdqLiLj0Vcd1RukBhvRPRTe0
uP+zp/5jq654t+n3qYowm4BJLtt64mZ3D4ycSPVLfN41U65BABwM7xBthqh8zLSr
R2KBTs1rR9yj4DCcWPo3a18hJzgSqseBD2vxP4Te+ECkrTRGY80LkqTpK5lR3wJ7
DHc883Vf6eiXpjGLdmBCq/i5qdJJCLmUVTyLxwayevyn41UKunPuvA7//8XtlZND
SnpiwTdON+vPA0phvpetWpAO/pHscxtNSerhelWJNsF0OR7vnBgSLHHEIrCYKE1J
vOb/LYYT1VCNGk29U5Ma3GTwJ6a548ZjjPkNxO0w7j7e39/dLByLYgcnwxX9JufF
Iu+GafYEXCjPBZd+UZz85UfeiKR2ljZ4CHC+6aI5xhufs93SwpE3Zw/usszq8Qrs
8se1yX5/AZ6RlH7YGQwvh0ct/pNgzgcTHLd7RGaXXPukylPlrn/iQIxUQK8dlrCW
kmYqZePVoT/Y7x/bC3m7sugWsMbOrvRQmwYbmL7OaPsGlGLjz5tuKI8+hZ5go57E
zeUL6jeeqBOiQ9LwEQuzdYPbkvMWNNY9eR2itRhKelmdLz4h4XPSfXuvtH5t7a9h
ioQtmg9wFg2/TaxKXpuR1v1klN8w+aUA6z8dbt7gk3LowTDlRmpmFvbUrxWmp8GI
2uCSSJpzam67iYhTraDiInkzAGcrdl9bvVDLlHJwlWmsCt8wFMgXeDnmZvL0TSCV
9erE8S+0LtU8P+7WsF6KN1zh1EbkWLQpkJZUOrES+e2euENg0BjYUyRV/aSs0msI
gpIIvuJVF3pjNLzuMAwy7lPbGsakW0R5+LFiRYkeI20HvvyhZDHDzqNpgXGVhkSM
iBRX0t94OFMu63SrWWZhLk0x5okLfT/5J1pc+YrWoDuO5wyqp0n5ZoJ2fBaqPoit
qAtG8LDhyY7w2WkhoMTB9oAFRifnWw/97H8isauKxXPH8+49DDvTc1s+AE2uLLic
T7wx1seWoOkEl1mAZ48neUldfQuyTLGmmr5CEf0gfIyjnMvGiJkH8JEzD4S60JrP
lpy6rjv/NZAN3P9snwdz9p7oVFxOONvJYD44hJWnOgbWlnxe4LJ+fli8st2SB8Dy
LeNqlhGFE1SeEfiKWaACQpj6Jc558dPMHYn/g6aclgtspVxH/MsItca31gjorsQN
3tQSdljhhTJA10TPXd6IBUWYfMWXF4eDp+JmCrULlMDK8fK9I8XlChW7YTxPGg/J
OahhA47rLqbX/i3hHLGRWLZ66tvEHmgkbOxmBNPiB/31my5Ibs0Lxlj9syULTaTX
25WxsG898sI6nX12n3jIQ38GW+g3ukoBPdbvV0RBFg8Ms+cDGNcJ+ndaIFTYx6BT
bgPEeGgNJzzh/SNf2wdi2USLb7KcowP6L8UEaUXUJUgR9KY4s3UH88D4q6DPGaXt
IcInnZaE//3UhqyZ8cY1Je4xWf5DHFBK28cuYHW8lZfRHtElMZasTZn9wdaUtTIa
WxEdsMv0XrMKGMUCogNzcxBwcv5xpu2nGikvsHbt4Ccg1jTalO2cH+AN5oRe3S2I
5xC1BeuV+bMhoy4n+MgEuhKhtR0g30LRjngkZvJvONrdXMRlJSAwL9kqBmTLLxnh
TL1qm43Wehtx5gbN7Ho9Gz+pGx1OwOFNhjCP1BwFvjfmjUvuSm4odsLFWW8xy3V/
yQi/PQwSbHv9EhZLFg4iRHVKvbTXQVAaKEbS4fKdBFwFG8NczH1nVZmrnbvDo8Aq
uD/qwOTpyDeXo+8kVda19AV9fsEYqfrhgKblCoG8pmB+xB1EmyppwD2XDMoKQjgM
FOkImfyJrnRlnJqM9SHpD1bBx5r0dxOK+H1tQxp0jSYJwe6CvrflbGy3FEI/Rots
c9S3xKaZ9KS8ueo0NdEzMoaO7mkfWaTeqHJG1cbTIqyBQSB243DbBQ8J538HT8eZ
cjgDyJy956ZLMfy9Jy8UkgFS91Uq/aC9sLvBZpXb9SAH3658eMfJlkfnqBAqNqqC
VRCyqaQCOm+G/lqf8rr1s35j3R4qupN9Om5B9r9zOVBiinhE9rxhojq6jQ6+tDeX
PGrWB1xMBtGQDTjafk+9nNj+t3aAR0mj7Es58VRTI0RPaBQRLOTCA+bQtYGDa8Qh
iRgGKUIlTA0DBa7PH9hzeKaxvZASrNOeZ4I+1ljkXm/2E7p0m0YZ3tkJYZw5khyZ
JxdX0lqLZ003Nfke4Vm4VEX1KIbOOrT71NA2PzTEjchp7HI/82J1eWBJ/nlMfExk
rU+ZYJYuzoeoCnbgS0RL2+CAjPdGJd/ifK8Znt7/8vNOdfp1sYwJeiMAYGLW4pOZ
bybFy15waBK5xJql/CA7E+9Cl/dBskl8xzJxuZ2n7mNIZXoi8SZx77nhqpR+wdVS
iz93x+KVZ+3yX2DP+uEP4RswOVHDIzJv6JFkzzT+BF4ogupd5l4e/qJ6oG45pP+5
RWhzf80W5LfIJiT4HOL3DYiZaXw4ps1OhHR+hwtIF15UCEY0I1Y5xzhVKLsCt4R1
9L9nkosM2x3jzDd0Evf3O9Vx0S1U1qn+uD+2cDWuDmVVEgVX82AJPqdUzGD3yUnU
qVygVycjgmar4of7xFPk1cxpFwOkHp8J2VIVmcScd+wAd9GWEFYbBQ+HbXgx9gZV
aqcR/yuxJo6nE+YqDrOcEuamnkOtTmjZdiQOVuo86Jdwt/KfBXzPj2Ce30eaDj5v
ZIWhIDkC8EkAoS5jkpCDNoWDOZOUv7lDAX7SGJG9oNr5ik7tM1SUGwlYEtAlyR0m
znoKpJfFpB70W/zTXoefoKW847SX2Ypy+lPDETKYl14CWkMyxcvreRiRYYJKoFJ8
rxnluPvazM8ep+bLBRDgI8goQcvTa/+HZKMAy3gf+JVOhQBFb6uWBbTZQWDF0dyP
yEKrPJPlEY9iyQPVEDlUzrdenH+NrJr+EEdmIQm6akgw8I+9tHB/UOqcdliIhxxx
WRLHyhffsxt/1TYhzHCs5Im6c4huaE7vD7mwQz2Zh1WDTsvaMF7jCft73gjfMXaP
mMEX9ODiG4GylRUxD5ak+cvCcqf9OBldWtRIlMi6OmWGmH09O/mSy1tCFu9frNy0
ribpI5WiYnXHn2nJjSVM4ra3X7wcsCzplCFyvCZi0I2DrSEz+PMWeUmi3UgA5GNq
julgAUvylYgzLDxQpt9uEeEJvypjj7MGd4vBj9oBPgaSEM/HvRo9qb0xiFLhPhAf
AlFbrmk7D0yC0T0vCtAoQ5sqSLGEgmKsphoDtAQxfv70lhQEa7t0+4THRyIXZo50
9WDuq4EENIhnZ3pRiCngroIAVkdIj7OPE2lAvLz+N4sytbI2G0W3/b3QYTcSnhJJ
TOZKhmThFJZerz7aymKyRYfoADzj94xw0jmmBs6U5ecJ3QRUajoTddG5e5FWGOzS
lXgFp0ukV6NxMwrPZ+5NLFLLR4xZxnHKSBFOC6JILpv/IDIp+nREelqBo58lts5v
jYqY0U3/lIbaY/yzjfh4e5NtTiEnSffgRsggS4XPuOojeMudaPLWmXQ3Kx+JVCfw
3riEZ+kaucNH19uzYGZOYNjq7HkAKQNJHrLws2DufLQH9c2/8GsoWCGm4XHh8JXp
2EPdm4NasBOFKr7E0X81s3LOc/tSKZ1cxDcJqyrzBZTZtOQ9BvU54mJQPqT4oV0X
zMeUratmw6ctM1vJRvTE/L6YzYHSeU5pdCwp+fKoO1MaVNLN9xToakOdv9XhSwzt
nIeVEd4hEavY6exUXc8ZX42mb3dS76s5Ibyy1x1uZBDfxV5HvJfZrIMaVZUVblMO
/ZvXUBftj7eAUCSLR2/s2wYg9C+xkakjIGuskwySLtnWoyx/zwiKzwRay+jetyvp
pEETatsHREsZZKFGJQCWolJePfKOyybMgLpR7Uvwb8E8QgC+RCzkvUfhE5EISKAf
7GRCNQE1oOK+o94wTL8HoQOlfXKZuqHszU0F2oyCRaK6MwE/3trcBgVeig5v4faQ
vjRA6sSD+gjIchp7bF4se0aA/agofKN54V4IctvVLTpG7vQuqguHkmm7/iBpWRxq
cK9KN+QvetpmCZIrb37SOXY1D5PkSsAflaNRwK8mJoLgRUV5Sl5vhrVrVQvOexmF
OCWyD+FFwAVGcyrU6e/yHSqpvlEqmR9YjiUQI5OZFKWg/Kgll5M5jLSWFS8w/Kdh
Sbru88J7Bh8JaxzNM8RSOD5aEwA2I+M4eBFajrTBUvbKw70s3brrWKRPx6J3jP0T
R7jsv1Nw2Wfx41HEOtBD0l8B0cr3ZuAoIDULCz3z1S31tXb/79h84Zy+xb0BFSsz
oNchgkTW5zfFFoEpWwvvMrU6rkYHrPF1Y0JrAtLMAPvrfodCURO+h4N3g6NsC/e+
9mf8F7XzeqbLCweOOYl167ShvnliCClpXBbQRf3arCVsAfr+jHLQR28DWu0poN55
octZhdTlAzEtmaD2KsBQn3QewzongHdb1QBBnmpnpkGZ2KSYeGOuvC6dtvGKcFKO
gWzHjFMIF3D0BCKMaAqmrBAPQzNVoaPWYw6OE9D92hyPRdE6I7cPkD2MweWKJNSZ
XBtzE7m35/u8B9xiSsg9jnL2HbYIZM93se8NoP2I5S+5Ylh5yyI74BPASrgKYDHR
N0+AovAnBAV/UjSulDP4TlJVFRantPCmnpvsdyTGVXXzswOJh0euA7bWf8qtYLq7
UMKwaI2V8QQB0Ogl85IirbACMBNKgPVWqXmlcr0dcEx5awT1PsTwgOVPbHTHTBMt
p5cNlV2cT9Ux/JPPMTJsm4/oqylfPeLsC2LYKbOda5BpJpjJ2EDA0APy1VL8bR2J
Qn5npas/z7AnzuuxX3JQ1XmQWq5GGMtPlC1rQqqq6O2M4DVt5yAI9uf1xKZ3ul2J
GSQxlJXqHlZNIwydc/IGITeOmGvWAqrqvz67j3ymG0vtxHnLC31UnvHHVYWYRq3n
iGjq65ZlKGELVzAWgVwlLybLoM1n1Z3yF0PLOXzADFEHcWk5lOH7NRN4bcc8fevK
giZwD4G1wDxE2WGKZR/E3od2Dd2cb3MlkEcAl47BtAroNh+JSjiVOKB49AhIqpGa
MLV+mpK4hcuUmMFycgwieXIagzGAGoUEXg+vGvsxTaqhxPEZM2FJz+yH130i1nZ4
+OeQ7SUlPPkZDaO5O6PGT5eAGx41SjtyUdmmd2K8wIq2LiYnv3OlcPipgMxP1W4s
zVmQkZ1Otu42nbzQA9HAgaM4Q/gnu7OzbrOFBPj9+ykKAEPO2W6+nTd7tUWt9m4N
FIVrQHcqcE+KN3pZ+wRgdYsZ8dCIExt44boE8z35toBd1woZBo2HP5/zxLz4iIfx
9//Zfgt14SG9X7LyePxe6ICeKuW9W7eGtvoaFlg8vfugu2vxkGCBKk11PxDmBO22
1GAKP1N5kpe+hdZUAaxOtf6AYr7Kl4ib2FeBWOjxNsNFFUWHLeUeGuuBgBECtrWR
1mXz7pwxRve5tSSW9iuzGA06ljnz+B2v7KvmwZr8c2F5NdO8QCj5ZG7emw1/sipT
4JQD0FNxWK5YvnuJG9g21VITRnNychL07eVYM8wF3xKCbOh0ZQvKYtSejIoSO8IB
5lKjx/IExNL+Tw2tUqBIqbLsqkJTiiLOVRTxCGIo89rC/MFjVFYt1s/cuKgMoTjd
JG05fQefh/G7l93vvTL7d2c1Ka69BEaKvuZpDh4s0rEL5uPTx1UZdyt+pBXr7JVw
a4+bjg0ipU6CNBh+TKHjKjSEF5MpnjKzJHNKF1+B9IDYiT6Vc0mjevdKFAlVBrBv
jw01KlqNOQzVeab8RYtXHSnN9gmB4PcEvtLFGxpf4INrZ1W9v0U7lJW0pc51m1C+
+RPpa163C+xGvlw4I8oWRevSOP/8OFrdj62jf1KL0Egp00ZilvAS3tr0sl/ztMkC
C77YszWo4XksEzCnQKiTo0iX+RGehgnBDt1Uv5/CDEUE1Snb6ZhP0Ft1VACcAzl1
TWNifS4mXeww70jp00Offtp/0qvRLXZZUFNZhW+WNw6w2AzCT4pot1crwaDt2bVw
Gbp8A5FTbJpq6iRoDFCBP0GIKCHfGcuG+XTDo+5IgN15Xf6nmgyhhJcHcXDfOmtn
i3caHlhhTWPrEDwxSLrP7/bYcn53cZ5vfWvJK3jCXFLvAS2Tv314edlpZBZa7GvX
xBgxDGAnIjuHO/jP8WArqo2RURHVqaaOL4DWW6zATj8Zq+h5RHD8BhHUJpNLby6o
IDEX/BDPGAq/rtp02l0WPERX4eWtPmrj/2yXrBOqfKu63Pfk8HVeDrb2GeJgxAKl
LwBgSalm39ExfXUGiGIwR+9HOGv7Lx0izWsY2LQR+NlsrDrMd+Eae9KZMxUtHlog
sCOPkD+jdfs1nT+uwj26jjXPOY4EAM31YrwV9THqaCm0GdCnaB/Z5czDNUUy6iNP
g/qpeny8TYfHTEXDvo4vciVwjP5wcyQHftjFl0l686mR55prK4L5Xq0BfRwVNXn8
dgHb6CF4PLDyPmcz7iNfjxWxvyVdgk9EVoGr7z02ivdNvoQJavXb/t74vXk+0nqE
cDksEoFTb8cBcO/YDvYBCoAoaiyr1c0fgg0Z60JTGKQm+GFszsNO7iKdFgHpMdsX
ToguyUcxeJNdnif8iDEnK4DVIuxEwuy/P28VQNfPSlsGs9Wo/giw+YDHmlhd+Yqp
WyJ+5Uw+KKTBgcaXLVp0AegMqEMfKFhrUjxBYva6+QYiSpyNKa+pjQUIUlsNkKLM
oqQ2su0r47rMtMfUur2qm+l9LF0qeJ/SUFic/uWj92L8C01GypbEKVVt0htnk08s
UG4rmKxWR+YWFLZTnMMX2v/GZUmrdNgk404tzEN/ESjStcPBR5CoEnXiDl2BaaUg
dKlQoPUqtwKl/u2JGrtj0Pk5UicY8DuYqAUx4CMW2SxcljNFSHa/YHcGYgl6wG6o
qn/jWVrTjtXceCk8ecI8GPUJhlaGYzz/WVdPdANlrfRFZ/LzbQwVerk6lFxhyFro
knHPdyx4ccRGh+EMuysf404WUmnYxmJi1qp8qR1qYuwWoWexfWCJ0sZSGQENyHp6
3CVgeNUAFWGqbq/Nhb938YzZlCPLlrmx7NIFy2ObVlWXh6bDmP0m1+2mGM5uduyx
NedGXbn++hkYPfeoISqjW3P6CcVYK+3QkBbKAfgSq48MCyTcCrQLeoZRk0Z5siHc
YAG3xeTbjLLMXZbB3zxnQUp9It2w2wkWuhKn1GxaG+irEvtPKMp3PlW6pmZD1Is8
oEcKxDbKxWD1hpwtMtyfaKbcWjHlUMeWcGa2XWYKSU8Loa/AvfYOhlDRooZuD+3H
+hWr03BW1dxSkS6vmysmbqIHURJ1gpp1QyGyoADewc9KkIzkblbCcK0yXuwLHpW8
8N0Z1f918qru3KsIZqNFmxMEBvmLt1db6LQhBqZ11ABGa06yjhqDcIeFlgFk7zpg
SR4W7YuThdAxMfNhDqfIFnPCucYnwdA8lyZj8ALaZiy4pl6yvFk7XPGv1U3iGXuF
kTPXsHZRhq+sM1sNvWyUJUfJfWOmR56wcDmTj7zziYlElaBCrpMug10oZTI35w0L
pu6CPLX6EgzUEdHiFqnHOq3+0Cp9aKDfbozO5H163z3Jt8lq8jgs/9Oyzwka8YkW
7LgiZosokbI2xFZO+33MhVvG4V6sEg3tFxY1bjmlm/+kMPHnSdcB65Bmnlc2SznZ
R7ZTCGZsBVckK97r+fzfooh8Cl1Maf19uD6jgqHPMC/vLTs/12d1E++a87m6R+jD
CR0lADq9bHfH9AbEzXJFTBOtpIxeBUz3S2g4nTrBiy9sk1k7KGiCBlB3cQSd1bI1
Adbr/ltrgIszqXKGeoe2aMCO+Ws2MGsPEt0FswHDQ1BxwHWF0LuIwPglSoHn6gqZ
zTybbta12dgiKwA10jArnU+irYBSsdcxcNioNaFiZDclqvMCXqVnI3C354fsC83c
smpaeZZeJr0ZUNBRcKAFxVq016tYVS7tDYfjsC71X8ur4B3Xzzw9ZNJ7qsp4Vfa3
rWhFaY49ulUfrgs5aFnQrXyheCW39Q0Ittp1wa9O7BMIPEIAjJq/IepDntzUbZpm
scOti+SBd8rCI1pcnR4OEqharZe3Yfmdn8W/b62xhYpTZPH7ownvrHav1xazbXKG
OC8cknBktIF3JsBFv7IWB5IiBxj7AAMmqwYOnWFwRatJaoJPrDkBHtTuCB8K8qUZ
vCFkMpghpOvoWbA32q/NgviWnkH68ZhOwO23rTfetPM1/f4tWBpfULeE489GsXMJ
uzSNsnkV9Si0ZMs2bK8GWsMMTl+ifcYvbIBr8O3wLQNohxxgzsYlkedRCfrNYC7S
eValrFSw7Dn3+pbjhOAbo6wHLOi2+WYgJJKClR/AyK7aMWQm5Z/hj1/C8Dczel+T
5foxaYDvFUU9wKqQP4C/0yOrpZDoNRbkamBZJvfHJqjhT1I3j70Jo8hR5uCKKhyG
ll8z7/dhI74eO7pe50pLr7RI6tdQsNahQXzXdOtypKB686GDpppmibiEXpoOehlG
3/AKgI5dgSs21ufOKI+7yzwgKuXvjnGhKuSitDPlRPXTiP2/8avmiLYQmsMVXNe9
vTu76gIjfk3B5phgL+zWliYdU+0HrS6p3Pout8usATKymv7ktlIaR73S849hmjGn
4BLN1okp5KNDlp4gSGI7fOwyLBnI0/JodJ+SnTW9rahPhOd7+I6LGea676oViBR6
28fxPAWu2E0Xn2XzoKA0rhJEhQXkKq+D9WNmZlY0bHPTl9kKupGRyQ0cPx4uaV+m
1IJUNESJac1eH0/XlTt68tQfV2hACPMgEk/U7ZukTFbNUYSCHIskBtTcGJJSCaCH
ICMIUgOhAk1rvIQIdWEnfjTz4YYyk/+T2QiQBYBf0MWJRFWlYxi4dH/fwlhZxwYe
IV311Dz0Xs+8sgOXbCS8pB3RJ/k97PCiT8CTEy1EjWcuVRNcvI6Ai9os7h+R1rDW
QjRBcVWVhGDt6F/J6NR4IMbhzfKKrYOVHQ0DlK7GkMNK1tV+6/LzBg0ceQsGXfrc
vI5BqAC7e4mEwFDCy6XJqwDyHf/tGk3hm26YUGh0vC8Qf8w2vo2bxx2yu2DWiThO
y3rt7H6L9XDzrNf6fEAnDcL6Yzvj5VEw/psSu2kgedHyNpYh+OC/0k3kpPu0yl/W
ar0ZZKmDN+Cm3GBGyULwcYiDS/p1rwR2ELRc/LyXUCS/wKzSIv1t1iLvw87tOiR9
GpFqHhY11Sd5c162nyqGt8l4Mcn43e/2JOtIMYFsHZBoyByStGfZd+OMUrAQu3ej
UMQ7FFB94y6ENbDGmf2VniirCGxcjMjGjcdPJXySGIrf9XhDfrmyWbrtj5VBHjDz
DRH4Ew2E0kNGDwu1nF2CNFBnlHLZjWdk6fx9nmcEpwEWvLNQdbDMzyYaZ79USDTz
u+9Lww8S38/bLpf+3WxxFaWNL//Med2mNbVwPJKWF1tLpcUrq03ZDvIwPKKb/F2I
Ttj6SeX3z7qSQ1yvF9nrT96hKZzX/QriUX4YJbQricL+tpRiUuYWNzB37uSY2RHk
UIIJvQwdRarO3w0LTzlwO+mJzV9VUJVrBIO/RRWlUSZ1fJcc1HPSOSTbGOoLR6+V
aD3ZWSrqgAIETJjfjRDz9xtz0lyZlPKQFSqQJkiGh0nSHgRzhgG2qY4DWtLc3YF1
yOenL2K8ghfB9oIGD9pGZx8zYG02Pg8uQ8yBXVzY+IsnzjQOD+zKy2jmKWMUema1
8RoXqeAvXnMKqml3VMChHwGosSzIwl0weuvgKkfGcz/mItuMN97tnM7/H/boOD4f
n5M/ESYONS+YxJKVvpFLi2tS1np4R4NEdRdvTiwmfH5GzTiT3gyUYV/vV1vqAhvh
Z64czND8SpiqQIwEpitxUKIYx3xv0QsbBN3bYG8QDMfRUWXcBVIqjJD8PsioEIDw
4p+iaI115EIxOd14SBXWsO1H/uggrcrI6WCfgq8eOM9VbW1eEwtu14rz0u+atce8
SLSBjOmJNkCPkolOwRQ6JiQr4KV6UX5etE3W/kZCMKJO9+DE0+t8QMBzzJvQLJNl
OyUMhsf25sd7n7dJbc1VA/Rjkdh+fWWlJWwZN6pEuoYBjTZk10xjsiEQJL9KluD/
cWb/7XI2rJAzoNzq2sTyFbb5oSfODKClRAu4YvlJUT6yxLPScq7nRVYv2sXAI7MM
/qfvFI4ZLjIJYGw4wMB+8YfK6hkh73FPiPCha7D1c+dU9FCKRoOoZ4wdNJGgIKVi
3lams0cv97Bc2ldM3iu2Ua62o95FbiEYN6yuTfm0fVVf/akE9Hbt+xuErNEvsdgz
rXOLcxIR1qQ/fRI/Kbkbv/NdrSGQgLadSD2axyqRYf/ob+CcqgoIdB4vZrNYD3T9
CdJ+JNGmqncQ6MzsWEuDtBJa5wtH3pV/AaBGKtp3RHuWCQrHQqu1mZq/1VDyyZO+
/DHjQ1AfniwLDe2WthKIuD4ZkgqMRkIp32aoVdEiilZGb9+ZedH0Wlt8ezGZxHvc
iCpAw/2Vb+ugNNiQnpHhnmDZ6s22xqcH1NL/HSalRi9BKgBJOs9/wo/ejz+0PIdV
hm1DqoOOguQyUy/5jCVGnEqOy+qVAPnb44qdr7ko1w7lnc51BemRbQzhezRTWevU
7YjCyD2uBU/GNxtbsDtAO9j0IdSjjXgJJm3SFAGLcObHYpQaDa+/YW+6TsQVmumw
NPMhwuhMXBWqndm4a+ER4wqfptGFCxfNom6MVr0JzW+IVktcBmZ6/5WmdfuX+rVL
/KKNiXU24Oxkgd/Qs/oJwq6xSJRv5AgfX3AE58NQSXxpJSUXg+g6WcTapSn4ET+6
oA8MUv0Ea+EkHcqJd3Uv/SXL3RL1Q1i4x8zXyRfNXumFZHFiz5dMwEPk2ILDCZ9P
6p6rbknvU29+PkmIIwo7ylg8wGjp4jMa0T7GG1yw6S0J8rovluXcQdOBgbKGXT2V
/YCUGtqH3tNgzdvzdBaYLRPhmXm/IQH2FZJPByd3AI/ukMAAteyVJraulwEssMQO
Otcb1UNC8UIY96S5n5Sysxb7+fb+sc04ZHb0SAA6sBFqlCyaqQP2WkE9+CvLCelK
HJtmOMSI2Ym8/VJ9GWiyXDIkTld/rq455SCsseTWPncM5p5aPiNStqMLlNevmUB5
BUHbjWtGrWpgKIR0yN27VcNwODswJlVS3HPKrExTA9K3dAxu54NayANq1k0jeBV6
bR6pADzFNWdCVc+Ut/9csIw6PwMUdhhIoikljMHDSOmzODSyhNtsqpwkzyaK9fze
kTJLhuCEVdh6GEEyqsr4NSMW3NR64uIy1LKiND1r1nCkQmnu+9Rtzb9MQ/vrT/ra
9hZSllNIcJWqTs2O5GwKRXrwrrWYxRwTQaCYdn2VofVtYtSPJFJnb3GSiDpxsaiY
1gqZ0JGr1zlD/wThU5sXntLkTrVywDhaCnQ4JVaD0ujGecgjjzjgjhhfVcNRaFKz
whlrfDRJFrjMskEu/vxfDIXb9D5qW3QQtVMh41IiJEACILvyNC95yjQIE3HaW94Z
y1J9dJEIzqgwSSSp1eKslOHvdHkCMSHCjiq2UbdZrcLLnu+tsmFD9K0Ec4270WI1
mqL+6v6ugbVLkMrtuLY0hwfCQgLOCnMjZEo7Bcz/TMQkHYrSehkFPSMWYqmrNIU8
vh9b4HFThoW7Ju7dMU8fO8VitYWxEL56FCwhgnwUv6XGT4nAbmEZ11eaUfFh6wav
MsQPlPCWigl942bqPxuI5lG1k0jUTgR846yol4iBzJoDTlKoApVeLU0dFRvzd4g5
oIrWfZPQTPHnaxn0psboGG2G9sOrY+Tr+TQCQjybicK3I+Ugfe2OJPeR3zPofb9G
y+nJq5YqvgWI4aJoftrYtd7QjuNyNHQaUf2gqm4KlmI0jro0z/VP8+q2u9pyO+gP
Man1h4TAR0tAia+N1L5nck1rhgpXIK8Vr4ml9HyZWhgeoT1Oz3DEz8IRdt0E2WGr
jqmWJ5qsRPpLNm8ht1y/FlUWeDTckJfbS1jO/MV41lmZ6aNvGR9Y6LzUvNPEQkCp
WUYXnjNbJW4LyDntGtNxqWJu3PYS8IHTa1icnW3UwpsKL1oymfLuwuA0oBwKKdRL
ncjnfRPfpechyLvLeLFy+zFRwGCsVgYwgJ8Tf5upf0R6LZTM4XyOjueSsV3Rf/Ce
3WEGk2xjXaTMt3AX4hUnMKglQon31nihopJJjCkozOskzWOzxx21iBBbmS2sHN39
8S9hRn896azii3WaWi3FkTCQlepNo+Fsq1eniIstOYHR8sMC6kjDT9xCjN8r6bgM
vR+rJI3Zo4gynVjpx3tMqSNQZhYxPxC1WPo35H3uXH8wAHPxIx8Ql7RnZNAGkNEp
3s3UdEQg4ky6UyBPl7reZ0OGw2qVYhu7LqVlT/qGhlZrI8uwnmaXrlWliFYELqDf
nXoALdUmALzmPfVi3TRnlcUB3EKW62QNqjmFdEvYA0M3MuiMTltsUq/PLDykB+MS
3NTwALmsiRuX/aAXCJtELrkldIpmEREbIsrvDpLvXwKlWukvyaLWqGunMV/J7Zzm
D166gUs3XK+baIdOhK8vTUJx6UpBLzedyKahGej06eCD4cL46hWG+Ha4cemb95TG
Pzk7DmFzsSZYwlZaIEBWP8vZ/iAFhwj3cXqlnI8n8fAoJA0Bn1BqDTQ3DxCtG8OW
R5dEt91zh1goL797oS/LTqOf/OPs9ujupOff7aq8gI5pXOfturwR7lmMzrITs/9j
5W5YEhrxQgVrPHuPEgPDNr/J/EEiP1Dq75CGXs7C+xIhsQ8MESAqIZMgKi2vvWIs
gy98mwGuonN/raG2ArANPX7bYlFluPzKBK6PWRP3yN4D8d2b569WgtpOT9n+SxZI
8GQg2YtyCCIHqlCWui5ICM7ogwJXqTjjyHRtnqi7qYUUJzaaCZpHP4u22sG3gMeq
EwsD/YRhOSWu1tkaSectYOpOz0T5U7L5zy3lebe00dSm5ZbTMMi5wltSIP/lpbul
M39mqM+R9I+gqjNUcYwWsJ1IjTySOOcQsD53ZGXDufkTEP73EVRelvEVNY2DNOGt
4eqGvjNaWshaqHzYvdEXzFMs03/1xbPPtkQKJNB3a4NRZ4ozWi74Oe+n0FOZIXH5
aQWme//rRLmVX4klpldfFzQu1xmM1smCMFygZSINYwobbE6Qqs9DquWokhzxibZ7
P5ijAYixmJQsg+iww0X5UZvTCvnRCWRIN0o6lqVXYrh7YnTYVK+f9FsmB0qHRvQ0
Sc2adPOlXu89mYFvAkKohURFRgfrIl9IkJ9NMrv90K1gJWLFzq57quV0brOHzCkt
/uoE2v85QUWGeTC1xX7h+2MP7w5sqJt8jqCD5u122JlzzoUWw48zacDjtUxx8B75
h/kL7AsmSabrIIAc7KNq89cRWWR0EYvOd/0H7a1KlrRVyjz0CetJL3q4TL/QDxaw
3z7jGOngKUJJcjTq5NkweqZaBroPv4AyIYZ3F/lkfhHqY1z1c4KAnFwkbzbG7dER
P3VcTTzmQ4CFzza8GwYwgwghjuTjWh4CDc1iq5ONPZsV7sEaQpURWio/vxNAP+Gl
6lfqFftmHhR9IfMWtGOW0HmDucO6psdY40+VSKDiZJkq9NqXfyUNgV0OayCBWF68
U+FtMar7Z3Y2MvE7EJQHA3FpG/v4LhxvO6xwiY8qcZ5d2QkdihwQ2yZw0FYh+q1b
gvBpJUv75FhAXXfqa7o7M+cj5zGBbDPCiuNtrykno7/KxRFVm53H/8UUcs0lzStl
/pYjiJOlTuzbeJ1NRVUD8IHbXRIwFtFYc+520xmSN87ugX3Ps3p4kSa/VZWPfgCw
Hmb5So4Lr961ve4YMSGPHYh69snH3Wt7wf/8tB+SjqG2pBd1xBFp64QmZWlGFaJl
lWROsRkJGsKwy09RBnLMlokEb2ZQRPpLoqmILsTCtgnPaO0md5vnbfOu/nOr4PLz
2fJf+9BTUUJLz3dGkoU07AbFn5/2bpkWCrmrymbcE8udx8IewRQW0/31Hp7CnYo0
zYJbfYiLFH5lOcyVSsJ6KVlvGy8dRNATo5zODcgCOPPM1NrrH1Q3OJmCw2xaosxh
nLhQRgGbKensmHqMOxeOhoxfhwQayWd6p/EkFEG+CYI3KuQL8yaBMMkfad7CYv1W
g0i2R6twWwe+d4Ui5HazufT8VqyGH5sj10bDfD8zvuh7s6dEkuhyAsATFp+h9MBY
drBdeAH4k6w7z/6qwNhscPk+a17WCFcDZyrQ+ofEeG9MTJ3sKNrT/lQZXWY1KLjN
CX5+br/ooLdSI8l0/IbCxVAakdo8DZ7pvyBZLR/VRoIj4JYaMczf1eI72bVt+26r
eJDGvW4hm3r2062SGlP2PlcRxEWThdwrK7K9pGRw3iUcUc1itjyVXzezC7rtymGZ
hlgc8sROnr6leIbbVoaPt3MrOMROoFbFVUzBbQ9zPKocbUZyXo3kKfJAzsFWjQ+g
8uk9A3aBIYXswETJJg4pRdbr4L62bUTR/GnINeBL+y5SbGh806wUqIciHyzMouDD
Hk0VjTmPd9DvIOuWSARPTaPR+vXOXwK2e06wLmo4NUUp6ZI6toXKMdlVgRCiaxer
DjgnMk7DV7IbAUaHA28otI1/IESZd2ehBJPOMQtXPe0ahMWwUaiw3Y+xYdjs4BoZ
BRZp5rw0/GLMkZ+CFO3HmeXYEai5dFOBL/JamLYIDDt/DVcQfDTN3+UiFJwKTXvt
CNaGhxUdpZzedvZLUahLoOA3U3iywPBGAuGgMp3nNd8Azc2IS1qqYHHNTNmWcG7R
ehTgNdjKESPuHIiNBfS/7uYbG2JDYIEoTFloCKqEQGvOWdyQTqvKwevFYZGX+Lkj
HxoYjaaV+HQTsn8+rDldqe8mk9e9rB1MRq1osJiP61lmI9REXUcf1Q50Mhfu8JFD
5kXgNUvfJS1HCPZcNUmMVN374UaFutSRvmNEgaoCVOuEY9CbQhjahzFfru8FbVIu
4AcqxBS+igUp0J9sqOwAW4HwonhKlnC/8exa3zhu/rzUircE9TMBiYf2eh9+ylfK
xRZOEwMnIH/r7cApKCHFAzI1VQGJHU55VIQvXEy6Hxbm8bDs30Eqk8fO8UkkkRNR
HsvB8FAyqy1E6FHWXQVY9gYcmfNUobCWrVZYwsIg6mimjZ16e0GmjihSLbaBOY4E
nFoSJTXgFgCKaUScmmvHl3jODcHsynuJ6wIboneQytMSdc0Aq5fGLSFg7Ii+h4rc
+Y18FOrvpF7sWKLJdvUragG6W02w3qWVuxdmoAFn3cMqAQQf2KXDTsTgyT5LRmX0
9cyjztAN9sfSRHzN2c+Drm614eIkNtjN5dz1vJVP6gHkPqFvcEDzOZ0lY0ajRfC7
s9uPS+xLxHRCLT6V4wV7NMC1Lp4qteoZN7Ag3LimkJiyjLlnbiWVEGfn1Tl9eCUq
zcSNlQA2baOQM5PnTyElUdjYaNT2o0uvy04h5PmwqRfv76ZFZmCMVooKYUsBiH3Q
EKFTKE3NICKzQ7A+ED62CDwuh6nHZuFvsSkik6M5XGGOeOTGC13w0YEPVoovxLYu
4OYd45kxDvNIbS0U4U/ksAnzEe40Zy1Xe9tyL1mvw/PJYedYG7x5ST2uLqPO0l4H
cDa/g2QaEmsZYHjKkdhd7RYM/dRAESZXk4KAHsaSHMmqKNSejligkihYbnDcMFuL
2tqC8hymqDTaMihCRj3kLy+5yK9wJ5XO350O97y8tRBga+WauqSxaE49pjbQWoMV
Owb0299mPuXfDylIsPrN1H+BtHhN3kp4p6P0EzO2gzZ/X/ZRv+ijNQ7G86WcFtIb
uLnDQvpiSZUAsHHmTd0RBUZ/emYz1pJ9zWbccQX2cotyTHkDirU0ttSiJD4Yixxy
KIQzoByzms8lpsiV2zQCNVIxyIgIMZf5W1daPEbZNvvxUrCPqA9gSyDNu4OVD/y0
Jq0TDPhB1lni/J82r0PE+nrUmGkMxwdAlRn+QUzZljz5UHsgM8snYUREIXkFzR5k
UeHirSp1usiD9AkwVXO5TltyTk4rt15j3YBEPy6GTrfs1Qn7Jpcj+fB1GaKODhUv
gKt0/bbdaFUQnKT35yIrQvhR6IDm8AOcecVcgBvhDFBD5O8WSdEy9hktjh0NGH8w
v3bp2eyUhWzVJNY0r6DcYtr2LtShEwbpZ1oRLFgGuaivWbTFuE2QteoLgp/ooSuf
shoscaroBsQU9sCmh+5WwFF/+kmjUH7SR7mvyqaDpmvA05DGKEYlirR1Ayv2YaEr
yKgw+k/eHi92tcOwtnJ7ZtuHYYOssErys0SfduvO8wTKXD2prkVvqLKB99iYfoOJ
Ul9tUxJh6X4+s7ZEMxw+/XFdD+ICdXyoLYMrfaAYAUn+wUSaryNIsRuvi9Lf2sPJ
Qg+CcbL/+CHWKMu8mmismgCGyfbciWi7Hxoh/DcFJzMXWS0ZrjniHE7OcBJJAy43
lGjGbYxnH6JoMVr8Xoe4QfS9DzXZHPy6t+O3PQ5H0owuZJ08qqFRdrFa90L0TcOn
m8hgJhyQQ6c9+z2r+sal1DZDM9mEfMbOqRgCFTeJg9lfuXVCwfdiAfmXAXgBynBs
3YXcMKXL8OtQ8joDDuz7ajrgkMhdlf6Vxj/L7NiJB8TSeAFjwxG9gLgRJ+G5UCku
YuQRofKs8pZvK0XJCiq1B7473w1EONaQYcYa6ftsqqia3oLcOWQS5zWdL35/9VMW
S0edeUooZ/dL5iAwVcPJRY9A6U6qSs4CUQVizy2ioMr7Y9O5SaCmIM5s2ux+8YRR
G3hWAfLSZbkxfMXdXG1BUW7yAk3j5HzBhwKs/ujXKby3y4z1DcP4Hk16kDQVIvBY
WRmMTXVFfZsJQAwr9y3xfzTxC1bHlwVsxnR01XmCIiZ8wY4s5xHW39R2Kn7l4krZ
OoOhbFYNigFXD+nVKExgf3qzMjMm0J2LdlgvIZD2uKseSntJu9DfLpEYw8cO+Uys
p/t42Z9GGz0/14yvq8TVOms4SDEM6v3WCH5ROeJv2mjMhM0Y3qI42Z4RrxDfBXtX
7c7vZEPS0NxODxG39XKusdhXdfVudEelYITD/OsaX6QrKjX+DvlbI+oj24OcfXaX
Ii5KRcyXMQu7FMohYF0zHNbpJUZaIsh9DCfis6ixfOA6pVd8Yf4rgj44sKsVj4oD
Crosa1kR1kpCp8dMRo+zCXOwiJjYXNvFKEV51JU2+dD2B41BZ44Bc/F9tVWu0N7q
zpoL2ZNkrarjBh+t35IoAvhl0Rqw3jQNnool3mhPPQUyKlhXTCM1l8GR4HwsUSON
Mt+aR3qGA2zfh983O3ms0/VIZRksVzPwxVXw7jv9dYv9b7l6ct7KpBECHJjsy204
oSvtWhYyugOg5akMupSELDPwmRpjE8ZnQHaGiGOK/3v5UX+COUNL1kp1+LNt16Tt
DXnJNTQpK6pO+8VgN8g0foI4jxisuY4213CUcYZPgDC8K8Rn59QwlJfXBzC6xxNR
cntyIUV+sJfsWjP4bUevcQ6/58fplEPke6RvhEuCb8b9eD7Ozzw78whyZisyuMEq
BhJSnUJZ5CSY9UtAhFlnQiiwaBhQrXj2YjoqHVWihElKsDiOeZo8oXKNgh2cXapI
111HG81zSpgQVrwON3AwPwnVKsAZPHJo7wYMzHbBxGldxI5rV85v5qZGJ3xDS8wG
PqGaVhHomo6K8erEjD4drXRsG1ElxaP8I6rTPanR7datnoCVBWePdcRyfApQokhs
PBmTcTNADv5lvpeESj0sR9zm6+A2jP86y7VNKVi/AIIdb7TFDdeGzOFpMvYa2V/b
U9/WwduZh/Loe7QUHgiB16ubDtjE+QGGhnxSSBfNBl7AANxbNe9WLI6tVS8owpx4
91n9c0+VE1ZXVzFUd7d6YNYiWNH1T0AkJlcYIt+2E8BsR055M3FKzy0wNQQ2mpBc
5UNCFVTYdDPn/a1Epyr1d5li7AY0TSxvNU7qK1uuLIIt6pUxd+Jtg5TBbr+AVTed
9RHVToCyD2PASmqmW6ce/fBSzryBXiqydTJz/3kJRZPBvtlnuDBStfvEWi7W5SGL
vaY26MlusvAgE5CEXAj9nrDxC1mji0r5X+Zbi7J68SMV1Nc4eR4bIcfcnKw438Or
0BmlDo2hNBR/dg7VQsxeVX3Tds50Kc9KBHH2ZDPWo5fjJGh23IYvk3Fv54xQhLVU
XipY55gQr9S/ct9y5Gy1tCINMf5ebaOhE9jiffv+EM82eiUGk0rnJHMr5AHveBWf
b/wRMOE8nskmDcA9G5QqgqbnTv0Uz7nXX5NwSNGCaVb2jAydP+OW8166+GwMERmh
MTQgzkoPnR0eMK1qo+BANctqXj5qlzP8VGZiOXqF80GNkAzq+Cj4YfITmsjUFYcz
GyRbZh+6dPTJTgFTiFxGppElxEgN7ixOHyeTalZr3ICsiE/8PSeW/NvLOzEMWReA
Eg1UzhRI2Wfq1oLUfJSJxxaeOcU87xqcR+pOvtC4uwqbsMtPjLESFaH4duWULn4w
Ig6q5QaTx//8B1s/vNy0A/b+T7HtYalzOxpMn1y9l32Cywswi9a66fBtxTsmZJ9F
6C0OFF6KNdOA5xT0HT2ZliMIHYscTLsYH8J0SrdeOPLhnNf4iZJ1cxomyp+XGC5S
N/ZXATJ4xlpz5pP48L2glj9GRW7fsbnAkNogG0pchMTzQevdYZSN3PDw3CUPnwcw
ynYYKTtPge/Fe2j1wyj4qwG3kz/waz4rjix9rQOAiWqhd3mXDcjC00RiIbOJeuwL
/eBMZRF0tkG7nePwhoEexm/Y2nFlTNlE/RKYKpNqhA4KyAeDCLqzogJzWmjZzDbT
IyuG/MNaiGsgfd3wotx5CLxxsRxtE4mXklRFZpnFhGdZ8MBq5pHYAbnoQNMqgKfg
i8bTP0aZ2l1HJgyHLxJfz3qn/Fu7Gky7WU8Kr9SYcVhHScY5q0d25Af409YeH16Z
FmfCGEG4W+P0tV4NyEnapKV11LasSeAX7xX+yPDb2uh8B/iy4ruB0p1LZGCw1TGL
Sajw5l77Od/xxSb02Ob9Rpf67L3gf2EfUBE7rh43iJY62yWjnDu+Vxze53d5ftqU
uQJuhz4iiR80lNggNdwMzoSIVszvTU9YgO+b8/or5EkEYN0sokSCg0sgQi+FxUsg
v6vSnsXU3ZUzneCVE/b8KXTL7HUuyZPNKBjCSKSLN0OpF9x4bCvoJNlWNMhcX1AI
Uk2oMUOKenqRWhoFQH+pMqnnByFwpIwD7QWX3eeujYTvJVPjVrKNiDrL9sT8hz9+
TYTJjKYOxeze9ApsZZHHiFKpqLwD4QOfnURFa6xnVtDDlgoq4ztFmoLQ/UlHur6n
vBWzgnMMwJDrn4Inra9LOLp6tdXJTmd9grn0URSeRKKsWuxxJRvBUnWIqvWQYH6c
IPtF39zCCXf85AACjrLkSiLWU0s98zKBntGfiXleTsAmxxWiaEiM+vIWOo1wK72v
DEpVHkdnRO3ZU3jfuzsZSF1dug0wrcUEhbw2kZJTNUonQuB+YnQmZ4eD75YEA/+t
C7hpwQODgIi33Om38dbWIcJ4wq6gujV8oOXV1rBDLjGpjhSYkLEfQm4rkY7xpt9K
Ab1kl62vp6K35WSMcVyS0vWS3mu5pM2kC5R4dti8xr0hdsZPvREaSFOanzMWlOjb
XRs+M4XTzu35MiJHD7nXW80yF93wK1J3OynIrMm8DJUNF2u6d6KhZvuxP2b0DLam
5pFI2xEMznfqTxV6IGL86MlgjpyWxlL8IJ4q0SwIxs+wKzwBSsZHwXLDVRWJHfxp
BoCOcmfDBvRfqOGjHWK+BTSShx68f7xcYiNDzCaOymuyNjaVywW4K5hGR0f5Tq3C
NczmFGUrxZUElT/jpdDOaA+MN26A8aMtFYTaXn8vJPJCGr4ZqLmrbmadsqW3mg1M
XXvZZXZwDpKmg8JWgR9fXEdMFr9zdLAIBOlG9O4RJ6cgTIHvjgPVoj5ipquzU3Dt
c3PgI7IlPsH+fEU11dwT+zheYYCbh0sSduEO7j6f2tP65aa7xMGDYOqrtH8W7p6R
YmBgAIyobJ4F4xmO6gp5fWmhRPRTSdMGZSyWcQkv85aZ6LCFpTBkUukXRH58HK52
0u+R98SPe17jHrkAEwgpAEGnoqhORrx40AS2ful9GQIZWg/TP6Fb4icDLuAD8NG+
5PquguOYhO712bTD+FKX01VsbL8bqI8vRyqq4xyne1tj9UOK3Qb3YUwhfbwQfv6w
MuqfWWRFF9IwmhtGaIht5mpGLj8T+WGahV+Dvmczt49keLYkVWG4mu0RFk89kcK0
PgyvXPJpJ8kJfTfMXPn2Hl0JTRdWxwJ3iQTiprOE1DYo288XhyvFho3UYA5ytoce
7lsf8m/CMUZ4puTH1aNI0+H2U80nQO2L0+/U66/CIr5n5bxiuzKavXy2r1vAhPiS
F3s3WaLymlyA+372ov2SZDy0jJUE8Xfw2eJ51cg+quyq4crZtWdwQjZBT0W0f7Nx
L6QX9D8o1Mk5dJTgKLmojhsUFSE2ojFzUvZr86R248FlQZWa1xl61logxquzIxg7
fDyTKeDADDah1GmA1DiqgvRs5FBJOxi6ym78D4Osx//B/hpyv+ve9wj7/W4Jbweu
z0oTV3d0fz/3o7bKMWaZneXqRrl6cAIpdB0DWoFlhoIxe0Pvcij+E3DMlI5SFHUT
/K9PfrgA9CB5i+ULpieAMSFS71jYMdr+quMK6PUHJq7l5iYQCXHHcwJ8UOgHT2CE
PNUZJ9HMirx7e/4ukWSo7V0k19PpI5iJgGptBVHoV24or88HOvfoHkTbzwvfdtE+
PxGzvXm2iE7RBJ7p24e34T5s46k30RiybRAr8bSrx24gyp5R0V/zIKUKhBmfIKLt
Ux7FsshfKRhEDUUxYW6CYzqysNVzzniKXce781ihW8e8PzWgQZPNn07Ln6Xr31sW
uwmxuemmuG9+0alMie//+W2nYlz/fMQux+HrjKA0tIOcf2JCjhC7zXSbIjlufyou
4JR4dlbILFr2CXl7+VAYqhxqN606y8GtaK8pMfjVisERVIdR/wNTve5VjC2WIYZi
sOG6xU0XaPtf65lkbME060lNgRoZDFS6A5gL/SPO7LR0UXj5QuR6gLWEBDllwkmL
zXhZqLIQSspxfzZNX3dfCyRizhDCVwABvdvKPQyAWo/WdSAbaVCkXRyw61GV3W+U
4mDiE4sYktsSocx+j6t2cpiHVdk9GLHqrmWFvb7Sqzbg1cLdDuuB+Ou0HodxsUyZ
xqa7NRT+f/idvr5KZI3/5pEae+16p39rgLqFv8AB+JxNggUp8k2yQlnvo+Eh94fd
dk/yYKvNOjkqezOhVEu/rERJJ+POGGsk2CI/bYjAupJYShkPAUXxUdGi3Pco/YRZ
TViNviIr36g50bYStqYrS8BziVbQ/SSCFMoPcu9LVj6D4EcBAlTCC9s+gRhhoEPi
3O15T1akrsavImU+X/qyBRFFQkM5bOqzZvzkV1ZQrgzaCWLbOW59UQybE6g+mQhA
IQ9Ntm9q3saNVE2WtwmYTxdigguSNJj7hVJjIds2jglrBXceNXfZSDDCRlOz24t+
nYRxU9UqP3JGW2D1V0EZ8/1en4kWnxM9mh8gIS28xrpJ6jSAsm5b1CkEU0Jm0vyd
QDk1cSo7n1x8PYK3qMv/q74Xt+wPuUer2FrrgpVNuVcPmlJQXMWNMK+bBxXtkpOY
geD9PH5A7W82EtbBHsZoM7zkQzhauamjFGrmde85YXUL2CXDGd74uNrAV+QBia4G
PaRB/qhw6+Zn5d4wiBdCXRpEW+ShDYRA2l89rLs9hIWdmvL1zE8NqDjCj1cOcIAA
ypT8ZHhRRiiuExQVSGp3NB9822DBow9MBRjyyvs3poLJfXE5SK3JDNjbqPwTuhVT
/hLFfBCAebIJF+zMf+HseOrZioHuWTWV0zvpIJSzVn6HecnM9SBUVX7IbjvlviEu
qWoxarZvrxmv9H27EumKl08Fpndik/GnHD8eWal8Y5Y5GHOsujeMyOFtRWDPjGnG
3A++c4fISJNg+JVQ7FJAh6a0BCl1XCQVCGQx7LBebGg38UlWJ2WKWpyTuf2PfHA+
yvWh8rzSZ5XWCM8vYUM7z7Xh/4ODsnLG0oAxp5Sh7czfo6SpMekBBbTcl9hrSPVh
y2rxsWNcf3tZsYNcrtskFn+2DeFCIyTB4R0DJguTZHIBoVPi3cFkKgbu803qWqBJ
qaG/VOE4ln3WNiV97ep60qPmdBMN7/jZIk6i0wZhcxSrgajnejJoaUyJlD8mRKvy
P7DHLsREIicEQ2uT0dmO23/Vwp6aFduoUUxJp9Tx4366OkpJ33ZQic0CetktRbw8
qxnwLiiQQ+McydnmThs7mk0kyayQ+b7WrZo2PaqV4N0eCjW3ovwPOyKzUGXaKGxI
DCLKUm9dYIwV71bPQBu7UXVait8CTcSKD1kAUb8S9uS8e4O8dsSxzIec/QEO1qFk
1jgMYkFO5VDN+TWHHhiPhYgXPrx2qPGoog4UvuiRoENkpPZfHgHyflrZ08aF2bdW
LumwgTcRDcg2RNqs3SGEwTiau9g3dU5O9qyhzrqc9BcnVS6IkzFb/mQJmYpwl09U
vKzhILOcOOzOAklvnqR7iQCht2g+XeuQX8xvRgwPamJT3DEsbriiToJpdI4zCe3j
gKdFo5M6ZukzwyBOg2OjpoGJOj4+XjKbeFDoHMNEI5oLofaPQFGmRH3dBHB7Wb0V
zyEgjT5n0AikZeaBA8wT0F26pafH45fL7ZvgZwFLF4igXUenW8A7AdnrmQQFwNI+
PgUWSAJZp82fxN1syxldVdlBtk1cNX+b38OdK4JniQZh/5DCNwtPrJ9T0uth8yCl
xa6sTnCiEBkO9qt8ZiQEI9a16lNuUV/z0UxJy0SbsxGjc1NvmJzHezKvHp6LXndW
2b5fP1JOkShRU1mMPCNzPEwQMH/6dePgigZDtFepK+PHnN5ETIY47I3AJI0+7/D3
dWEwdfJOn12DxnpwJppfckJ4AJJOSprOZhNSoykFDPmJ3qPXpBhaTYW/uMIl5auf
E9x6Hiwjup02HCYj5vDgXCqt+5tHp2dUVI1Pevtt5x+3ABpr+BCEqQzz1xPuJKu3
DCYTf2kCNXN9KDR/mzwyBiVHbuZSxEr6jIA6uPZWc0xBJn9CvXF+1XW6JAlVf39W
pPURZW0TC2N3e/0peBIOemODZauazj24zJoMZ+vCxh/K0Yo9ppv/rQ0U9vWeiUGV
5nXNoJ9O8vdJyafWnzH3P4K77RTn4jAFTALYBSCbuo5JPwFCT0+yg505umZjmgwL
sYEpH3IbVQd6epo3A5sNcgOIPHLWxJJLRMBBCnfI4B0+MV/t41rOkTEi1cv0AfqH
aNcEWzUQh0en5QElOPk9FfJ5S4mheGPcNm/zY5+Mx4Ww0Z0ija/YpUblrNPHf7kC
AU7MByLPrEXuymSKgNfFs2J1ae1F0R25n3TP4r40+hnrfW4hQYRpD2KFZq6j5lqN
VeR67/T6YHmlI2EQJUMjhn3IniA2U7lO6aRIEaNbgMCOlc3mEX5hu1FpgZ0yop/X
vEhNwIej/0IV+GVqd3hnYc+dEQ4t5ngYZybZ+cxQs/Jx/QdR5Oh+nk4b9AekEo1a
5itDlJSWKW76Xepkc88qWXAYK5WacvAAslA1zyU9hqG9Z+OGUSDpUR2INhylTGU0
qLoXvQE76uxtnQ3Xa4u5tMlCpTiUDVWIDsVH25gV/GINxhICXLMrsd14flcMy6MA
EfhlzHFPA6SRz4MGCHI77qOxN5TQAiT2iSmaNnhPs5GWHZH0ufSb7r+ZDNeetdAU
0ERoKCiUKOZPZRPxWj40dsqPhjSa70LN2Pww4+7T6WaAHCWaOb0BitBBtUtf+nzx
lzMqE2U2jo2dpupNnapP7b97ULm5Fr9q4S7sy1L2XO1jpY+EN3JMcBcL2LC1RTtb
oNMWgm0thwxdeoS6Ebr1Frvx6bzIoihIWiQqzLo9cPukfUgqvPcF5eJOcqa41IBn
WQwh9PhEIuaAtOSLNjuOqmd3NM+sqbKvjVlGofoNfG73Nry0gJvCPfo0pCBeAyR3
/Jp3AtS+fqIKwo3fcwt3Kv3Lvu4M3hwpmi9RojiOf8Sq5ANJbPyx1hCLyG5GTxx7
4cmXKnwRtV4GJaUzwD9OfwsxvOw85rut5NH0Xm2yxGJKTRIaQ5E0NAJHESLAlrCU
Mf8VyM5nW4gRkh9k8Pz22NTimBbxAU149WaDw734DxpJZxJjt9yhFnTcn64+1ITO
dX1dOS7WHPp4qDxNpS9HU0Aj3jMWStTTIGpHVPWzCULrsu6od5WozV8qQHF3wDuM
cn4J0PxSMuaTVOYV5af0xhRWAtvpXe4MKZVpi1LREBZ+rInhLU9LehhLE0LFeyIC
mXVXyMT19RIaB8H4NgNlXLuRkN9z3f4M64U7d7fjdzJ0gKUJV6F81U3VPS6D8ttF
FeD0VCmgL2dw5ynVQxjxl6n5sWThlXSVJV/WT4dMjMrrEW27d943xws22g06UNXN
pu4E9r3CSAuydvrQtJFrd6+QLEKpUYvAURhdrbpL774/ehqEy4FFgHu0Vll/YG9E
LojBkUe8e7JYCjiZ7bwwGN/6+9E1cmzTlg0D+dBERLUZUREN4T2Hr3HCvjeL9kcS
WPauKbtF4GW7yOhRl7Pd5Zx/BxFiLwbefPrhxz1wT3im0KsxfTyXNx9cY10WpJAk
SZ/4w6QuciRoJBRjv79Li56a1H0giRySMtMc1rkir/gDO29uFSoxVzuZUL+av4Zy
k6663XLhUIg9HU0rOGrr7wrNA/hpOHvEGeTdgw+DEUAXRJKfgSBTLn3qaN/A9hk/
2mnWLvpogqxqEBqM6X7n9UMx7TFu4Sx4WjdtKQK2mqdE+/hAcRF2qchT/NJCdMZF
YTL/WjTMglgxpdhLoqHkUQvv0O/B9TJyNeCKllMX2x/ncBuB3egJ+CarN1p1cdvg
mJLTGOjVuDZWQuN6mT7wYIshtibHb0e5d2YGTyIxzBU2wwUYPEao+LLC5x2To0QW
ZVMUFDeBnO2Q3voZYWT7/ycqak21sqG7iKVZU8gJCOIxRrvvdzMoLUNkc6vUMMH2
7q/dxHn0FA2W/acyRV5XBuUuoky7+j6W9+/u/WOHARVynjrBhbGVb65Zk/1yC5hB
ZWPfBnFwKwobRu3nrco4uewB4ZFKPlPjLsCTEEPNz6zeFjUBqpLZgSC7zrv0uf3B
qnxgO9rhEe/yFHuus/QhMcJztggHuxd9YhZLvfKP+g/YjkHPRZb4mK5wIoeQn1qO
xwrY8j5duJ/mwvSl87GqzaxiZ0cbX1ueBQX6B5WlsiTi+G/pvSdD4MwwtqTeo87e
LXHy2qJm4B391Lsqb50meDoa31GBNcTKKuJq8VEIcmsAjdCo1qs1a2i4ELrzoNv0
lqHsniO3suiqBk/gYyrSZ7W6k3xMeFvHooHcW8x7l9TtKbEoMicMdTu3fOAUJSBt
/Gqk2v6fW/6Odcl19kVcawl1UYBsn4CbMceKJcn8Lakbx9+7LYpZYW1c04EGsBHG
/vKVeQS+TG7X+gVoGF59pqrQJ5eaOHvENBSJULsvP9KsGfWdAtcUI7xGhQTANcQW
s5KjtNuozg1gcxypPqzQ3Lzdt6XlVHNRBdqfwJ4O+yqcpB1UtkeYjyHsBaFG3w1j
lAKzOoefQ4SKw1xNI/xI1/DlfbPxLnd96AV37ZSWomBnMve5Wk0WHGgh5cq5K++o
Nap42uIm7M5bpLt0avhwKoMt0+L/dcz9RDkeYK3GlXJVFJYckLPNvyUObC3CFyS/
akY1lNuVOmJkNZRc0hLw68xGx45QCmxRpiPPw85XktW3zBhVa7dAa8i6Lb2xmAjF
7EsPu4ZDbLx7tnsfD/9e5XWugXaxwknf4HnkfL8PXANMNdB8OxYTZ5vR1n4z2cI6
AjFG4NFKz2QyZg3lTzyueLrTHb0TVOR16fTM41c0Yp3v9pQp9OLNnovwaQgj/ujX
xYlBnnUWOXbm5ubGpcwikTYfGFe6wzqbfSs5MmVFr1Bn5OA+9LcmAEYzOZk7Qlza
2A0M/Ku1sqCuwFZdg4m7AgO+I/bDGnXLwwnpFE0NVjDovhkbddUGLLtRSFGE4YuC
0Ye0vl2YeS26IRYL0B0qwtfw+9SB441lJp1idQOjah2DF11LfKi9bjV5WQV4rz7E
L3rFP4QND6kIMnhQLLnyCuFvGKztCegc5ETE2uI9nO0kPi9+oCPSfLbpMCY6bNYF
3JxGB50gU0EaIUs8JPcXAXpBXkCfs2D7aM3kI066jaB8MC6kKLWgEYXKRrag6PN7
g4QT9I4iwrpPwt9Jov5PQye8kNOyQD45lwD8WJbjRsCUs3huvXkRLYtXnFtUzxJP
QyWAtZlocdbHkw3/8GqnFn4niNzzN89fbUHuWn4DSScSuTdpXJ8sE9hHBp8A5Sj7
Myfbp0t50HDc8E5jCkj9K28ws9/YnaYeK1z/MCPnY3ROOvpKTBLji8o9EOkuvqXl
m+h5WOED77AtA5K9ywCTxT5tvjGErIXVG+uuKl8VoyyCWOIpVArJ6gkdka59ivwC
B/QHAmy3iptTizLmNl9/4WAfd/2jY5DOhK6//0ckreMMqsunp/UWyh1qZYy6ArKA
R7JVx3v7BZgic0LGNjWvd7d75w5vAohfTe7bIUr5BuO+x04gHx75gE7uNmW0TD2t
buS6EDvo1gBFsikyJtTYCAOCVgXzQhRbMS2v6ppIZ/9zrwAtEd6WGV9TnxchwMSl
///6EBM/qaJDsncxgKCSVYMgkft4RapPQZH1JIJlqQ8pi6A44LAAQiwomczH86kT
nBTeytoVCRQj5lpqPquIlO0gA76EwfjOKp8+LAlMvZLa665USzvoOXrSuc7Da7sS
h2RNcIVbIe9N0UY8TEGQ3G12sXj0cXbrXJpUVZkenZIJeIFT5O7s+EQsj8jzX5Nb
4IJDsMVCkawCeMeUEjkXQDgY4D2qQbCqDNAGIcSQgZb2+f9gLphS0me18kmNXAA1
OFWdKAcAH2B4P3R1cQ0MftwLg9oQsiTP5wSsrS3fRSPbXAzDy9ecQsUFmG6v60E0
5KPLVCK/Q1YzAKR8KRw28fI0o0VRZkdKMiUSUG3tFLW1cnAlri4KSQJ2VRm/rzZH
W30ULVNGcN4KKR2OzyjGXRJ8bHJyDrGxs28Y51sCsbv3sMDgvBShuyfcr4vqyatQ
PVffNbEu+vMxJ3rrSYBmCqRfO7coztJ92PEel2p14k2LomL25CR1OzAjqb8RYOnq
eLV0jlMlzQgxcd1K22IPDAFTxmRtFUvVyYYptZmClU6NpL1RXWCrHcC1rZ7NFlzL
3zftCnYlGvyyDB5FhNhXJQ8tuL1JYbXfqyOQITqgr+ZYeDc903KwbLLrVzHYFDjU
l4Tn4qB1t8oiR4Y7o8F90XeT7lpZRhbfGmQYfflOwlLLc6DEMIsF5xSpWsQ9Ve6D
AvaJpY1JQEZTrUxvYnhcJcK7+G8hM1BfH2U9bImQUuzPrRofb14UFdxHicru4Eg4
Yhd3ntLsCIAJUFhESWwLIR/NuGowVlRXvojG/pDqcBhBjGlUDSW0t4t0z62LW5Sx
TVCWLljY56arp0UY5DZU9K40GKPcAFNn3u//ua9IJcv9SnGeGrN/xtOqHbRNPKzc
MvVpvBU0ukcsjZfsAhmMMEregvkjJBfCf8RR/iveAzCTtAG3ZM5hJBWSmmU4phts
xQ4ymlxLChqPtA2UqI1D/XrKo7t1wUasb49hT4a28JwQw5jKSFBnd9CBgOZtaxn9
bibdzuMaznM4f9z4/GpJRSfZZZsk1+LkPCryN/xa/+pJxTUfn5HDuxpKtlyanMu3
cTG+6DIUg9TTloN0/AOFGlEGOgtQgIjzOrPiciomMM9SIlVryuY6YB5dzpdy2J5x
716iMBAWyq+915cnHcdYuxUF/awg/HdYf6WkRDLB7RUXt3+2ms50iX7aOFRZJuuE
LEARLNMVCWQ3c1wXHaobvyo8ai6oahIln0391n2npNnpnqOYgPBVHc8easedEUUc
vXmp/EbI9xHs2EFcsFzZkG4IeHKEzU3znKjkXm0Ue6zAnDDKWwbi+zY/Jjnu+5ev
cHFXVqKylcTeXgTAkq1N4LgUaVz8KSL+YWN0HhRHJoLRcCzuGwXJ5C34JEff5Chx
sv23qxPC/gKAxhzQq93qXBrcEeXmtilFoQ3lWAyeFz6mBC8Pka/a9QrmEiIMU5CL
05s2QGdcFMGwcrHA6mpGcawPUeYpbvXQosncS8Z3ubvTHxmyh5yJ64Xx+M3LyeAQ
xOjpeVolTWCf96S8mcfXjue5xLDqsqgU7NNQHPTkLjddAG+/gXua5TTBB7MdxSg+
2Gjw0EQ8PBwrzGuJX2LfxmSuXQS/EiT6qenbRUal41XlIOb0ghm6q9aLrirqTpLg
EVR/+95J9PMTvQ/JFDykB5r2wcRWTGzB0CTnDg/TVBlw7n3YlgEtJGlIv7/kfcgk
qIk7lSvu5utdVTUkshlINFbpVA1GtZY560mgOEkhdGZwGjgjJb4CKpnHj3Nolj1Z
sLrb6H+LLAgncgiwlVmg/omJnPGFU3113Q/qGucZSzEiLK50KgDIV5fLG4efT6OZ
GQO/3QGl5QQnLcVhvIyXjmlSeGyKKtZZgU3qXgsCcnVe3sI5i6Bjfd0sK+ckKlqT
ar7HH5OD+MLlxK4WDuSNiiHLs2VEF6wn31OxXo41TIww8VThJe/JZqiz7etEZnZZ
I2QHxm4uSzRwHpCYxvjTx9WvveIdhs3gI+VHXtW1ruftlzV/aETBz/oqixzSVcCb
WsY5dVyApEcqo2oGU8EHTHC5cZEjYsbxjJg0EIRelZhRg34y+sx9PUE3DpHdDW9w
oETkx+wMvYb0Iub95QMopGPvvOY0lMPE1vY8oENBSKrpqROf8bOVSZckJlDKCH/s
vSiMUNM1z0BUmKX1yILeFWatRW6W/GaJR8iozwgZkODfurA+kab8wAPB9epcEYxN
FxMh/EBom5pN/X/qORA8DrN2iU+CsK+XxFKpSiqUiocZtis/GxNHt0vGGKmeIw5d
AZNyVzt6+P4mQyF+Olk07FWHTIOHDS6JlvDF9x8xPmqMArndzLpMnN+0VkuRffUc
iZAJJFj1nD3UXOV6YobbuLQpTf5pJCivl/wpoPQB+DTLd2zvX2orAoudiWgGyVys
x5CPk6S7gvu88yarryUX6i6L41Q5kMJ69zc0wAHESXQ7TmGIttjAsmEDsnu1MsE6
znYRKTgwBXEZ/0iE5UOk577IJio/h/gtpSNg4lO0oOP2h17j2tnHcBpI/O+LrD/P
aVAUlepNEer6z6xkf7hrWF68ErwH1gFyadhe14s3v1BngLJmNdJjlmH1euqH68K4
aQTvcSfQ/cAl63HfFSZwCATBsqLbWK0Di/H9dMAyQeXIS1bYgZ+7CEiIhy4p/J13
rzGLmiEUhQ/ZUkwrKJyz7PcIfg8KOD2NPajfbAbpE9J2dFcR+BCHe+omm/UzO8Iu
gt3M8LGmO9sU3i1muhHO9cJUXg6yctaM4uU+X4NvogUjiLO9vLuyVcEo8ga7mDx8
IXf+LlgO0B5hOgYHJ5fXKkY5oJMYeJ8epD9wYrYDC/2IiAInwuJ8w62Tr4Nk0eLf
6ks13rDPBaFnY8RnkkjJ3RZaVNdhBfDvo8z9/DOUqOLnNVtOnPLNZN1JXSRSj1PX
qp+C6mug+ftZFk5R3pthb+fmbe4XuC0pPrAitgqs4R3WLRPMLmA/r1EcLjQ6fWH7
ulD6v05PaorxBLYYz2Q8gwHuG9aornuDaxbsQNpL7csIWZMceOTQZbMmX7yFOeky
x78ZUOHe1bp/Rh3WN2Vo00KuMuyTZYC6KAu9jkFOgH64nVZHnO6d0iAucxIYvBf8
+oHB7kJQWqICkalMQib0pZnZZO6pUH6URwhrNUKfTsc8cVkrUHt6rsdezLAAc4Li
AhPH9aa1oMcRBnDR6tYM1BDk0G4uR98c/gcKDsNlmBrkOUX2gfxg09pmQN6+BLEo
5QLszP2n/muE9ihnV2HVhNq/g0ILl1PbdqojM/lcwcmA4z508MRejLKkeBhCn6Da
3YyD0/7ytF71DLG81tN66T7Dexcjn/n4L67xszT4/gF3fKPCDc/QTsE2jtlvCFvR
HaPd5IlrOt+Rv5fbjPfeE57WJ1SpHBCkQDgjL6VmpB3XSMrDTIiuTz62CK4pVbOS
AmKl4qdLON6YAPoWbe3fVojylbmVXs4jesyfIjVv3mpFji6w+Ow9oasnHmi1TMgw
bg06K4R5LKTZ9eTWDExtzU9yCSOk8AWWq0ZGp0Ov+zGzwPYfLKiwFFciQ2RLVx0K
YxtJlSdUaUvffYtgpwyCYk0FlBPr651HlIH+5PMhdaysjK5TN28y3MnkNX482wc8
7CCyUaACOq+4Bz8Oj7q68i+hm4E7AUxCltVRBksDJDJY8RsS4mUYnwWCOJOnxRbH
h5gKKEXTN2j2VjZGx+6XWz6xKBQ+0jZZooacwca/clL3vMd42QIGCBqnp+FeboSN
2kKMvSpX3BA/ZjgBmh6JgK/sHEFEk5l7I6qr/UX47dN0Pca5u1vLDy4cTNsviZu5
yO+fJ7aIbDc9R+FvMar1dR9JSwTwn/mkqUbue3SaP2ecpvZWyD017rxInlHLq1Zv
DOL81x0nyWYIyIhQ5sB7qs8l+07J67nTvbmX/aAtx9STdQ+ywXfhGoBJWTwvLWDb
M+buzs+XcnOo8yqzufaCy7glQgUjRAV0xDSXwX0LDv/XoroO7zwFdts+F4/Xsl3V
D2t/AE7px93lye+PBINFtTRqpqfoivpW4DuxG8R0yn+EV/N40SXKmG0qwqtOaXCr
U8OaSUcn5OcFGG0YssbhEVgqecKpJR1lhgAmrTjiB8eIOtxDbtjzv5V9sFefwf60
Rs/U3tkBPxPuVL6hvvfeinuRhwHSHT1kumcdsKAvERwgNY2/kaakzWO8ocKu7aYF
uxsKEl3iR+b42yH01IsOeb/zwDKyPG/uaMEDcM8NkDo+0+Wn8ViFFfZefPJ8uxx8
9EtzTHoW6O1qoM6WorgVs4FNBHGTK0lGS+a34/zAUX7WDoM6v7Lq+f0ppl/k3Acm
pdVLhz7Be4Wkl2fkU/ST4GH7b30LtF8EanO5MT2wZU+bQX7q5BmaWGI3zjF4Pt6b
V0XCzjKr0Ai9hg8SGeOdbJR6iDccZvvj/Tni2iHxNQ7Lc7FIYyh2emKxNo0SkyDe
oguuB/Nb/3VK/f5anTae/YW9axrkXO4tXjZs4LrgkXLA9oPaj0RdVQMSq4trOhZl
3w614M1w+Pt81UrKXrmnuAWF2FpFD4J5tAueGdgAlfsR+AbxnSD3tmjiG5IAieok
Mlmj/Zhj6MwklRxtZkGHlanrZs3fnTnHNyZ7gG31fx1yiEtnNSnLtvCZMmFQQ6+U
1um5g9s/tiekFqkjS4Tsngtl6uLmabBgl4iIN/TaNnGNzQiivIhOUa7X6swZAsOw
KwhFbhDKzd6PB2BXIfTRZoCpmLqfqPu7gpdiEkBr4Nc9vjKF58TyxWhnslR8IdAt
rIJCje+5PPdP43ys7hYoEYhGUXFrf9hJQHaRE3TkEkQt38rlJTK2M2e0fvnkQASJ
vfjfStKYcRA8LW4OIMHzKTO2olgs/ToPRb/DAD966oIYo2v5Bxo2lqHE0ldRXkYS
49gImofStTrOjZavcl8y75J6+MpSTdyAiRB6rFHKwa30lHGH/bZAwpRLQ0yCnsnt
tuZL++lg9d8YZMPqlpe80dKO0P4Yxuz/KQPjwXrAZIP2SocG451fJH6Mbq9iXVT2
ljtG2thOt9tXWm5LuyundRViyieiIVIMbmnHPQ7GcuoyiCkGKIVuV7WwAaxMMCVP
FGIYTlKDamXRlIqLUm/Z+CZi+D/lCRmtlM5R6hyngZzEE2Z6Ivn96IBn3CoTLg8K
ZzUtPYQqMtLRTu8l63UwrwoSDHNNn02Yq9yfCrbOS5Oh/kXIipnaZfA0gakZf0uK
p79p5a3mdgUWGxsd8kqxk7kx/UjYSMyQpQer6U/3giK2H0TBqbIFoMK6fkDrnAjY
Stjqh5Z6kEXpjJd54OrMr8B8pW1pK2h8NGXAn9dzr1VZYvHLiO6xkbuK9MVX49Fl
YQTwB38uCCCFXeRGtUbHSonFjCMnEoGA5qh53WQFNcJJR/ynpKixzurCQyZTORrV
26f8P/x1p7MNT5OmWaSLYXWvJAouGHyCwHD5BWxb8BgAED9SaLeKIZuNWPmMfQp1
9BOYuUFpygWIk6fKiIytHIpvRLVy6+raeikm9vC1GIcA1x2irPyU0S3dAURYkGhv
ix/VKTUCZ1lrJJa7ZEknnF7HHbaDuNvcxJQFw68h8+tIUdCtIKjcQhSZ3GxzKhMB
PopyVBSud9KuB14ML22NsHW1fmagnGdbIsoi7Kw5Y4fGoXoN4o3pNICo1G9zUnwt
A433rLM+m9ToaxHVOBDidArwc3rfjCIWtL8o5iugOp5cPd8yeZfmAowKlc2MtChK
CsBe0BuWEUFvAUmA/bZ4hsC+TQO9B/4jtAd8j0jnSu3qftkzW7JfM4KPFD9lyB4F
rxtI7dR9j3g3n+EzW8byovLNhbGlSZtwDAjWW2cdNpI0B5lme6rtlFk4RVN6jSKa
sBMScRYve8jALgWsnNXjcHuwCKOv7p4AB8jmyd7tLoEFerhP2N/d5VoFN+ANt3Qg
0UdFNOSgsW9KNCzJPqvOtZrx5jAzcy1+MSNZs4L8DkQwoIe7rJepnUouWSbx1k42
TFSqoIgc8KYP1vq5t3w4arugZtr4JykQOXdZx2xjmDV7sJ8T6rN3x28o8IkTfurE
Od2IEvuXLLGXxjscPXu6ZE9Ct6XhaUivCX0E+BxhzAPTGCWxy+80OkICMaz4Qp96
5+wRVr2vnQSKXqq4u8+HjQs/jO+3iBqvtC4eVaZ4rGG47Hn6uffWJ6nhAxzuF7gZ
A91j7FeoApMFqHuFJYsXIUgmmtVhcckTGjRP4rqHBghMY7P0u1fBuwChTQEyVHnB
lF+fPi/qDKRlUqI2eE3ojmEeFViV04ztxAfLhSdCIzcy38tCRrHyxgz0HtOxJVKh
L1WUWlir6iaGiWggkZ5gSrQajefyuNXYIbWjMfQ+JGMU+QsD2MOiApkyPjhHYMPy
gRCiFodULy2Gi54La/A01XHMcYZrIrL5KxSU8Bi8th17K5Gw7j5jiREJYlNYjT7J
liLX8nKjINZLOeBsFW+XYiN7u8+ErEDnFa7ROPRnjHnUy4xfz4H62KDAENDo7VGB
FVAVMGh1IdRikndL89vMa4mOVPtO4zLJqUKjAE0NCGGlgKv7lGn5o2XKL2HZF5Y3
5726/piLo4gJ9TBJImCmKKIT0M64X/5k7NfRdg0jRiJrdrDjYuYxWlDkLw2/Le3c
ZkNpdxtpJF1po8jH3SvVh93FtyyedHn/Ky6JhgKpNx3Znw+lTVpOneXj8bHgad1Y
cuq+jyebAfkrWXfBM7fX1mV5bHV5t0qMqV70HDP6cL+XBd21R6Ielbt+d7LDw37b
qTcVYkwJZqUV79P7PadD0VRvdLIsttlq5VxfiUqo995Sl2grqPMHI5rS+nPedpIC
UNdhzjfOZoUmOcVlvGIofZfZ4ufax43Y5FbrU71cfvS31h37GxPl1/4hHlJKeQdm
b2Kc/wyshKRe8MX0uMgOJ+i53jJYFDBihVnnwfwMYosPyzWiSTOnWGTOMvatkDka
TM/gh6ikJmwTbW19rusmU0mE3eCiW9NPF74C8VbCH41fvl2iE55GvUfeVBfDpzhe
QLifOgTTaRCJGiefFg66xT5btmDifeSjRzkFF9M4zevD9L/lTkb3//afBY9ulsmw
g/dX2whoif+U61yZTVWYKiDTCh9f7N4UsoJxAtsrqEUZZYhE08sR6Mz8tX3ZxEjr
Gd7t5SDP56rrFUFojlPyjW/wmwj6nMIuakd9jKc+1fZsBm9tTVcqM5ABcKpRVFXw
Z++ionRzAmSBQ1eAHpHJHIW8Nra9qzHDJNny6fo8AP49Ua8+DSfLhoObF2MQufce
YSOaG2ZcmD6TOS0GKcEvOwHp24f59xLrWdaZ3bUOiZ6Xz+Abn8emJ7vfSSh6taJK
jyB1NyDWWUaXGGf4JOi5jo2fogYpKxFTZ15WU7sgxrbbevvRZZRZf/ZRiX9NvxoU
VAcBQaLV0VuImlanIUcvsFCY0mAHr1iBKnWd9MRF0aTK3h6fnpEKP/lx6BS4sMLh
K45qxquMvZpB+HPWvMEiB9gA3cpEFtCbAQ12yODm+5IND0HyxgMD+rSVGGfZdPf2
sUlwR1fxwXM46exmK/+PdXP3wI1eZGpTN0oRZzEED66XiHRqMkCDeVv3tKBWe4hu
Ge4SsAxBaaEDflEy9100jPw43Ip1Lz9o2mq+xOVOnUNBCnqs7Yci5c5Z/6z7X2q0
XiORo7xHf6iKSQLjaCth8/fWJ+UATB7qOsAt70+JqTSWguc8NdMrI8YXmT4XLdkG
0Zdg5r2OyatXPhAL0mtgP4Rx3HM34Sx88RVS9qWUKpTtX/SpJC7KmpCZcvdYXEvP
TIFJqXoCYbxVBFUNqdmdWvvuE/LQwmeanwBqg3P7PNiZHfb6VOHt+j6yfuHU+3g/
p3/oRlCkyAFVbV3DMzFfYmf7jtwhuEEU3m7khnsabpXyf1cyMOwbh+ApEF65zsT0
x6tg5S3zNJ9vS/1ay/E81cltDxzX53GfvSFk1V8NRp7O37fr1ExxSnTnEkX6bsdV
E7ggZ/73fpGbGc1Ym6SjQ7W3oACI63TX1l+WY3i5rREkRRFzaaKoM8dgTlTH3etc
BNneDhLOrTK/LmwD/YNSEv2/OpLjeeAWksmEEDoO/BA6pzetsy8QzCbVenDD7mmD
G2uKMeXvZdXCynOBW3d+jA2kwO/MtpxxJavxPbjD0DPsSaQBHnuXn9NOZs03jFOt
q2xndEwUBa0jOIg6oR5qMAnBBFgHe2U8h5k+pABVOhiEM4BXmdOAZLjBr7pvF5rB
WXnvwgALifIC26BT32kjJF4R5GxQoHH9ixvOLEvLLJIqtdIQ4VcbmiEUYrZnfneq
4itsBBth80r6Havvpj76EIkwUVDGx/FG05WqxuAC+a/Whf1nGpXha4KIziih0afr
x58v58jISJjuJyKIYOu2GPR+lbn8zw8wmIywNjtE8WZP+1ZGhwulBCk7qyjIHyAy
bvtkpBTGharOksroYdnlGMmFApqf+EpcoqIHq0//MI2xXi4VoXAZP3TMcpq3JXtW
0muQX7/WyroKRuaZVfYO1yQmzHalF9TGZw3tnaEf5xNFnq1NFqJ1YaNWb3u5PiGz
btBibDFgxEL86ZJWmpMmNC0u9zNY7W7K8u31iZgfqOj06sCjarbWU72FBsoz8F8v
BY107yE0F03tq0+ZJZUztIZl2fJMfCv0XIbZHm4rxCcAJ+ovtPwSGq8v7z4WeNSt
jx7zvZ6suj2hnsA4i/y2iDEU1WFp2mT0R49suhFgy3oR6vDci03tyCwdjMJE2LTN
yyVb8eeUBt6xatlBVJo5VQ4K2q3Yo+8es4ROOd+hdKLg2kGTON2KkpgqvkdAuRRI
5DKKv/pCSJtqHm+tsrIvbnIbJ2SXjMCVbEUNnUg7BN71H5k7V1db0WNt4asqpShR
kSD3trXD9G22KiyRDOwUUJ1CJZMPxW4/82BD+cwoLisvXSxOxQA9Em2UP34EFexw
YEr+f4BisDcCZ0RKj5qhgQ0vHWqK/bsibbQM7RMRI9TMqbqMX5Pxaad5sDVogVjF
pQqrENzP8ZLdx/7SE4boGFYCcoGYl+ClfA5cK31c305TFJmiHVoWajB7ZzoV1yCJ
+GYtz37F2pp4ViJLGKbhOp+stnAVSGzhrw4cNpP5oUB1/oa7ho+kreDhwb0rTAnj
N7n+UKlnIGlFgZQT8jmjeJ9MB94k+nr8DpgopI7HMJWYW/V75kkNfe81oS+TVaDE
Ox3OqlagluIIV+Dp7gvKJHpbEV5U5O/Q7E/rD9+Qz80yZOvoN2eTl2T1krPGfLVl
dpz9yFB8CyVYJ0A67lI36e48F5fbNxqtV9FoctsoqLiRYggqAXzxymq79jsMJp9r
zJw7X4uaJ1yrMJipkLCXCw736q7PxXTDzQBlvBdYCtG9Y3wtaofAkMhNn6MGdd4W
hxCcqCO2QxgiwW1rydbiu+yM2mDhcyWY6bX7BSuoqrCcLCYv5kEcXYG87qTx+gGD
jdhSkLbOdc/a4AHd+dj7atrcijLkNnqsgngcOdCc5WOhVY/9HVEuMAi7TbL6p+hB
yqBPssm763jx9KCkW/5H05nWSI96lE6UdTWygE7mT/Sx0DNeV8RXToMNxH0/3lnF
oQbQQn6DIPEDc/ARIkN9tPxTXoHuWL7Og8N85faoH+Gn5c94U5FHtjM/wk9QnidV
zvct4NLBYq6hUEC8lGisaUj0dpXXGUJhgmvJhBIytF09oCtPjUmAW8+i83X4NwOI
V0JeF8JkC4acnoQmWDcN2SGFDZi5xWWXmpK7WGa3qru3GqleqAZ0TNrXEEHzOqPV
SGrXt51FfFSErkoVlAZ+EVhPBW8TeyjW8ChnU5jkKxdDguuuHvZwf1PHBvMbTg7h
sxoJUvz8dZBuGQfcmMlcj2Jo1cHBQUBZsh9tdyPybS0f4gRtfjGk7wyMJLuPvenW
LqvR62g1xrKAbjuAmHQ/460955Xano8eKyhwjRI3vguOnCCz8wOYZqP2kgz03YgL
7QFniXjvsMYwctdb7xHGsimgQOyU687IXcuCpc95rY9y0f6SN1igNviz873k87kk
uLghko71kf6rlQRINkIdzBmTZ9HMNvDfThnNwB0k0DSVx46MiKa9VL2EJ8O+L43f
w1h4QJ1ka8/eiqtZS6Gpgz3LB65EmRk1F83SpK0UvGGbI8JM2R/iOut/RNKBap1v
wcxj6uad9f4IJlVpReCiSkBeaJxk/EyQA8LAGg9p/nFQ/yIOOgkPhwluJGHcAof3
dj2VfO82zJ7kT++gDyU0LJkRkA9DAwTlKms3I6YUEI1jZZzAx+LtZ7V8+GUGSThC
cMo/PT/0WVpP22SH2ZJVT9HT9Dz4TFxd2uM+H9fsxMaUc+WiPg8WeJMInFLYvQk7
toMARpJWBxw5xMKX/sd6efH5uE/dFiTmEIzfSqKoSJipOjbBwVKYWtHvJndBJ45r
mEgU8vyBivCbcExElO50T1zFFc6jkoRCbzLpURZE3nvlcsTJc8jNiJn69RFUPjoD
A4rBJFEzidapktPiasiJd91vPnr7gamLWK66w7IWhYyvjbzZ5EBsJTr2O3zaqFzw
abp01/3Ke0gie3Ww+3/eBt+KprLuCPIkgR/NHZ73pMIf6nttQ+Sh6GgL1JromwuU
ghoJBgpz/bWRUoRoYHJuT6px5HMme+FkBN72UrpiFgO47hl050QPBCUj7+pJITiS
gHvsfqcXbHIpX3vkGUJE9WkCuuk/gx/4cCYD7sNsthLQWQGqOlq2vwHwqONNMe3T
KgM6brQAObHsUfgU0Mfur0e5nNELoKJOezEuAGPptZLUpkggs1VNO0DWJy4VeaCs
Gu2xbfPqoBDJOa9V+f1Jf0h46H4NvPBZVUkLyCBio8QYpBWnoMAmXJLdE2BzqBzd
VSLa6E2X2ZODqtFmn4RM2rgi27VktKj7GQhNbCSJP4+m8EnnjborwRa07wzeUXi+
bOu6No8q4uzKdWbH0u3HomaMOpmDPqBgQ82SxnuXqSaoQVvBq+TgdiiE811WtHnz
bWcPwS2fWfUs9ZsRTBUETYeF8uwId3qgNwQ83/aec1wvxKQqBOT/QxNDIjeN5AVR
Erv5v9t+jmKW98L8rASNTJ6FiZhCHYGe4iHq40fHQiNJHvvocti9T24rklRmVnGC
2Is1hYEkCAhby3h5t5nLxowR89AOsnwiJf1Gb6zq8fGYlSrugZ71BVbF8+/CWiyV
uNaOlDF1M58NhNO9GRyl7Cy6jRjxjJoVtmBkRGZBplANkUxYrEinrmgDBWo7Gpwy
FQdza99ADYQ4P/Ydfh53m2x4VOyiBWR2OtHnb6PBKn4b1zI6l1zsVlsYiS4neilb
Nqs7+4ACAdKVDyFvYBa6LdMsSvtFcLVGNC1Hc70R7iAXdDZdq6PfXJfHaCizQSkA
/JD2IvqwM6hrEaGhas070+EkIMrVfO0AJsJ+e2xHJK3aru5g+9Q06bvJVhCsCHff
l7MfQ0pfGZH2owLD4LFRw5uia98kfvEF6N59fRREzHEg76kX5cvECOYOPaEmdKxa
FB8hP/b5hfSdMH8uzSiuNezirmaXB7xLD+b8OBWpE/Mc38K+i4BnxnTU/9ZznbrK
1l6sGCDk9fvkAZGR4oWZcTyxodPjpYHZGMLWPctH2V5XCmYZgcA7QslbLtdvVjGZ
wEDKuh7WyKeUf+qnobISfr5EC4rb0Q695o+HOuIZ6CSrwrktMo2/np5qNDJ31H0R
zSJ96YG/RcHSQHgeos5zayKCrwN4IUc3ZUnBv3h35pP7L4hs/WK0e0CLoXvUadSU
tjPVax9fcETCPA6s1nP8dPG9ZZyCIWcPCKh65yi14xfa1K/zJSsQvPdM/AlE2LGH
r5QPvQ9DawpNhFBeZ1nGY/Csqf0NZlq2olps3JnHN9k7CsfrM/dqA7ur/5b+k6RF
3bfY8Wpb/O8CmF+UV89S5U42hi3p9QwuLfbgvsYUjfih2CvxUShCpPy++i6ATOkO
ib3JjkckZ7L9mW1urzV6NMgXp+dWYCNOhG1mEFH+hujIhYqDqnZdPzwy7/nhsrNN
tiu6CEyAUPplBoqiHoMOHZF24bjAfma+0GXPOBkJ1io5BvOIvSUlQWJzh09kZw3X
+pOMtxQx3/0hG0QwLCiEC6s3obKZI6NMQJzRmkA6qtEJ3NXTq39HmmsRmRHqqLxU
U9oxW/EGn6oKG0bpYpCy3I5AptVym7MAX3Z1T0sP+EMG0B1yurGxtoK41tZQIhqu
W6Fn+BuPVIZ4XfmlrgYLBBrh/IT2/G8TAa0n2K/dxyiCL6yIsNF+dDLKSee1dTcP
ToXX5DNnwtQ8Gnh87CJyOIfQ2x+bhsraBON37Phu0VLSwwDrGrJkcf9t20Q9zmV/
4K8sJT7v6EcHx99Rgh1p4zmZTHJurJ5NU2ukyCBegUSYcXHTyeBxzVKeic/1S7yy
3Gu+A0wtBxqCHEERYGhAZfIZYw0Xsej2L97uB9AVK/QMxzdJuvunesZ9cxn0wdTv
XhgDFwiXeJBtpPmACD2eyI4WjFgmrA7y90KyOFdV/S9vB3iZ9YG/LT/A36MUSJCs
Mw1wMtQ3ujBvX0hnf6OXB0mp5VNFx44nEIYPaJNfi38gUrUCLWrIdMwDb0/wl/I/
6scqs7/sRYrcqrrI0BZi2h3k9grGqqdtcqYACuIj55MpEP4SYf3Kjb+kEX285/C2
zM9071NwLS+847G0/wYeb1FzzoQUWQnhc5EQoiQw+QiBnkrZbZ0ZGsViCbrH20yD
3LFkJwhOC4DIrw/ZQHP201ck4vs+5kxA44Vvv6zslydv0CX8tG3zRoJiE9Bprh6P
H2TEf1aOt6IGZEVsGJO2z2gOm6mxptNzZ35C9SDo17S52GWPDLEJ0cr0UUSJPhgi
uxPWQLCT9cykhn/N3O3PMtnX5/vM/8p3Q5AQhslAkBt9D3PAUEVBE+W3Q6gQIuID
SooWXM0m5UeWWEgUv8TNyRzVN2GZJqrKaT9Nj6pHwjZ3YaiLnhmf6O41lLRTehl7
OhRxhQxChuFSF9wwYFpeYWgo2EVLcuyFxjUX1Gg2XE6WzmnqK7JJ+Sv2slChbRzk
filJ0GCv9BsLAsCH7yx4XbP3e6TbeAnMGuIKbHmPoE7KH1AqWOzQOgZA/qjgSMIF
icKpWKRi+9MyPyft/NAcq8I5tfcNkZPs3d5cK6TfzURiaig4ij5ckE7z+PQWT+zD
HJtrNd+zgHoYnuv1VftEXQA519pI3w8lDPTwY/WbnfO/8LRTLTJK3vKX7dOzf0B0
nK2Jb1GG3ZW2EpkVlUcpiCkCj4uhaANh5GdRDt1Y+v9upmsVA6tj2Kg5/aJWnGXd
2ilpJNBh4VcPkS+vPyaASnHzsJ98WyZV+Bs+/TfPeUiL+TFZrN2aZsXbP88isgG2
Y00y3D2oJHdR5Zo9vvqtDxxgm3LW5NNc4Twp+u6oFW3Qm5I+WQJlaHQ5cQJg/MfC
AmOYmajBLvoAOLvm1f67dOBTIbfu4cIpN30f8fs9IXHbillWV/UHDAfyYy5DOkvr
lztHM4jFfJrKgZSp3jsSXtdZ4DmmoWdEhqgN2iHmDdFTzds0sJuY61J4FxRgg0xH
KXFQWb14HipUfqVv4uljXQfyxtV04G4O9oWLmKAuFjve6/GkbwG1Znpx+J57d3a2
S/bYWtnz29opO85QprMUjpc1PI/HNZsePOZmlisKyZM1WzPPQ2dLqyi9vP5j1eVq
oPyPkK+i0AKlopg6wLUgw+SThFZ+IlIkpXYLxNW889HnHDTNEufoXX3c4CNyfkwP
Z1tLKXSVFJkWccn7eWJnNoQBuLQ0wFEiBqXG8/amXsv4CzsfZ56q9RwS+VLo/nyA
j+EOuEp23xbDtmaot66vEBMfplOGzJdApsWS5wu7AptOSVN9OqzUcSnBc7tGuqxV
eMGQUlWkG2m+/LRIAiXsI7r5ZsDY3F9hgJeFTtvmbcBsyLzBdtKN3Zef68SSwmQp
Rj6MmnAStwybO8+AijLhHaMALOxaS24bYx12w5pDHYruEO/HWAYwPKHwByN7LLTM
dpgX6B37WW01PlZ+qF+ht71im00y4Pom2GfffxuLjf+nbn8qilTquw318Wvx9KtJ
TzOqqeRUU2Ac9cfDthDh/p8sESK66z4RC3gp6wpXmEwa9wFvtkoB+Qmw2cq4YMI9
OyeCuOMLTGHSJmRPdO2F70yapyNd2fsi8702s+bJz4Lk980JyARswuJLtQfiX/eH
aEbQWcKSt3p0PJNQa8M0sjRYKiXAgyVcCtVB3a3CRGDCZP8k44pnKERgEmuKDLdR
oDs1mWxfsv3pmOPcXJg5hh+jHZqRD9/t2Nse4XCn7UXrn1VeI4N32VJAX3+imxit
SN0L6hg4XRmx3kcKkI8590cBoBJPer9GjQV2FdNbGQdGUoJtPiHmljn5S8CyzaGE
aDiIH60o0C2hedczPWcoX6JHKiTN5YSWuyRv4lk4AvUWkJNMbPjpOvd8Kapr512w
wCDGjfuVnJ42AgZcHh9tMLpDY9rzenBIqOSOdpnFdxKMIiad6IBiPPnLfsMc+jiL
d5Rqszu39IJ2HjjcR6HLt6zsWHj9xV4hxQBpL/7g0RouYkIvDYEGt/o7kII5fcdF
22Rb18QNInD/Q0M7p0iN1A1rB1XXPQpQWGJjJV7xWxYFAQZ0591MBCXxYAMzFOMr
q7pggLNia2+1j3dFMkjuGFwNfCfaCib0ILiitlUsXSO/kV75J/hbSaaWiY7BP1Fr
Finx9connF+yvNF3SyHIVSPp/MbhbuChcSJ3lp+cyRFm/QSiw6hG/gEK4qMxmtoZ
6BQhjoqjbhDWBFArznnlaTFMKdoGlzsiX0NtP+Svxy2k4Yt16zvjpibMscLaMFKX
Br+TEzoJhgpVGWT5Z41w2kwRY7VnH465DKLI7qapMQPTzfCDNLRc8z9Up8Wdm8GB
Bfnl5GtCHcDipoC6dB+n9alHCJxa1d/ooSzoUnux+OK0F5anrPGINthOgmdgRBbX
Zio7GQN/ERfN8PU6jqz3foRElbVrAsSb+LyZAEII9zKWuHSneWx/IQB5J8j7ZMsz
oykG2JTUcUfgxFKxMx+rJR7lV32jz95O6/vkxLlo2xgsBAXl8J4MCCh5eCxoinzX
kluQiKJmFq3rOvfU0V6h/gtApRs7RbB7kgXh/3nCYRCySNZwaIKRtMQCikZL2tD5
UlX213NAua/3l/gZszSDuVC0ni7mKT9NDuOEcFDA2YuY5c1Q1CUuUmlsNjPHB4q5
TQgCo1WKyHGomT5Qa1wQLI0WD/g6B3Yag01OxhhMyp3Yw7MG0oFLDyVg96b3VREu
GmYdfEH36BnZgUnfYvCj1O6NtfMHSees1+WEHlsmkCVg1HtVygOGWEE3S3SsdfwJ
z/mnlzucqScTOm2AZvukv3W+SF/aNRIfOw8D5PZbxUJN5Z6JkDwBHMyPEdpjqNpw
7WriPlgMikWU54McgUHrOhPKWRj159uHTNlMYD1XEWrLnR2JgtO471yPxtB3vmPb
MU9FnFsBmyO2rTfkgUA+QeHbI9ny7/BGIk1sBVVzXViB1Y9ZQv0JahktVi7KX9pe
3GgngI08VXPf7godebjHaAgtYShGjY597g/sQGnuj7mWCaqtuMbhlj/niNF98JdM
6gz8xONDF0ya1Ito9BhxP5QkxUkOpz5M5NdYAn5tX1/q3AwQuQtVWpM63rfuIcJJ
zzAud86iyy6yn64bQN8+87XwDpDAZUzz6GuT+KLCAs30kc5bQhCakog/AauBz5lD
kgqrLnCUl8b/r5ET75eOYWbTAPRs0l78kSVKayBlIBWgwl+sRATUEUCdBAU82ATd
s8wGmidYG7TUzxgWkLBP6RWVJLOTxYfTvQEz/FLksw0qblueJOd+HenX+UK/sckH
y8x1KfGS+0zSmEsrGmdFmc/V4zmOznYsjieclq9KdE6RpqtMpmtMkJc3hnTupWlj
eHI4h2S9TG7tVFmz0F7eFstO9DgO6PbhwhC1mEBbluLfiDfL5EFI/79cArXYK8Pr
xinWmMAjyXm3V8WA3XJ+bXsRSxjsAsdEKhaYV1c1o+Qmd6xcWDkN2wFVodt6oczo
3qpe/zPEVGvgjjcCrdUMDm4MhLgJbYabQD1XL0OIz+gFzbTiptipKzD3XOvaxbKT
ZfpgB6XpZoqg41KfUbNzXy6ahfoVOj3e2Q8/3z0dOEmhQbJnVsTABogY0x10+Sf/
eK5UFP/HVTpiF0VD/yYkJFmcWpSY0aI95WGG90TbRJbGPGcgZC6tNfe1g3DhP+jk
XEqOTjt/Ic30LJitxR65mGhuZvUtMUB8FeyGMWGT3MtJdueWGrat+VXodrJSGDxp
rXB4xUKp8cEmMyYhvhaw2EVvfKe8Y3VXLUYRgPLRxlM/c1wMBicUwzBAPRTj8MsE
+Z7AdKBbwAyGpzhyBxjkLLS1t481ZeRmFM6S/88zXuH6/j5Hm+VQo8Dwv1HOUft3
gzN5f5bbkHGvY3AZ9pyw0tLM75Un80rCNDDatb5Gm5R7A7XQofQumrB6A59DFPqF
sfymgKyg3f1qDbK/n/Bx/rBgaF7lYGPQm8qFXLbQ0lGIBtLQjSa3ZrFOBPhFiCjj
RqHzpi0/QvnnMCVBaPonsRliW//CvolDOsIHOhG3Is+/iNThTxAx0QiFi89+huyE
umiDkyF4bQok0vb7HZLBZotj/mTIvuXJuM0ypyDZES9DXgJA0BC53OpcyJ3VqHgw
SMzc4yG6S5stXluX9MZAkF2V7tt21BvnxEmMB6/zWDi6d4zDm+UoTbP6r1PhGBK+
tMv6aygfdFR869L1uWgdjAgrW0Qrmjve23zVWQ6zqreKeeWVjduy4DjbJUM3LfKj
l053RbXE4G0g3RACODdTkGjvV+eTP+MyPYp6zvvqk4YnLcQmGlp0vy2PqupeeHUG
9mf1avlQqZyftQD+LT6VHJTz2dtKPYW7tJYuS0Zi/jndjmzc0ljutVdQxK51JCiO
sWCWppJizZV+ffBLuP1hdsKaLmxonMOXLWy544Cy9xea20/ix3letq+yyam/KDmi
Q7hfvhGwNCJEHlEpUnt8p5O7D5YjYmfIJTWDThAX5SUXFPw+GQh7GXofJDB/hP3X
hZwzbcAvjWKlrC8Hm42YlPTQtHxCzuimjU3o6y7X2akzHOzOKYVz+oWv/TA9657O
a3QQ9OBNbTu48WvBmK8hAItz8J77XqVdWyyAXObwdioke31jWmYhIPEs++8EgmMN
6vdytaKnGkRQh2m9deotss0nrrPwfLZgqtdTrq2Tie+MpUe3Fs3c6LZuRIy6U5do
7UMU0RVqcFDuBRnnFvQZXXq+5Crx6jskTVI4WWj52jowDPLO7pNaCmXhfaMXoO6j
KTErHN5x5keSKWGwRtkZQJ8xgFRknA53jwvQKAqYlZRmlMxEPEZhV8eRU82FaNfP
lp6HrC6dqsXYoCG+RmfFobh6xlu+uV6TDMMhWaGB750K2Btyc9p0Au+IRe5IWVq3
uEoBW8rn7RX/648H44BCEQpb9KuB+h2CjWsy6g6KizvyXtFvAOKrC44w1icCkxIS
aSEEQzEqHD6+M+xsgUxbl3CNPdUMWcxLmu7Dm2+7DvoC/3aoBM3e30CUDqimtLeQ
LUfUIs/sfVCS0T73nH5hwraMa2AgfgJRpeIizcbiGcaY5ASeJMOu6i1JOOTS+Xvh
ZHTkjDtKmuM1Spm0pnQ0bPFbfShNAVUMF8PnHqe5y/ARJHWwhga4PjVnb/MkpTEB
2BzId+mUXKpiy8JgaLkPoVh6fT4XqOpOV5pxDiU4I9AwxEvmXKA+xKx79HofCEel
a/gjhBqjIVwzE8lDJoEm4eNKtZY6VXcuSLTHbxYfusl03h2QX+uMm/24593mFtcw
qadoQb5hUoxpncS8k5OcwD3VJ31weaYLEavACdPDexRzD9pA+3a3EfqCJbTYkWCb
8Q1SGMe6+H4ndM2k12gTgTygPIZuI7ZfBO1S0bK0Cv0L1hbeZWPmkBl1QAQv5Ddm
MLLy8cQXWFTjXJ6ZtnUzmmpUAEtL2ruw2V1eDjOx0VByECFNDpdKkQI/4lpjGm0M
8anJ7WtG6refjc2WM9e2w+Zsu7cEIbuwdupHbNrxBR1+zyM25mUAUFjv975jpdrt
eoFK8rihlshDfOlckBS1ReQ+lUQcFY2bOM7rWOKXHl7n0xiqXUbfZVa5gDoRJxlP
ejGEc5+OJ2wzkt5moXVDTWrTqsFqTlEQBBqEp2UyYdkw9gCDOu/fVfa6DhJzFmOE
d1QoBjTnuz8RbUYLQmxkvAa+Mjq512YYPL7Z5eMUsEd/u7K4wSuLMbsqvKWuINkI
gsu8uw0q7jXfIfOXxNHA+vZhmFDF7B0oNUHJrVD6kx9t6nyGh9vWknjdlMVIchri
KS2d8YwToTeOd2jlO0Kc8NZTWcFml/eLZ2NQCJJrppowiyO76RFXHK86WiVQATlx
Zo8nZGtb0w5AePuCzKGRSNTs+//VsG6JXiRVPY86jxGhQM+zQSS/g2Pz9rN9bYSR
eF4tvTqjcKNsV7pPz2lJNgZkovOHrKGMCouTnzzXkORL+DffmlUuq8hrWNXVb7FR
0rd8+KFLT0yh0R/0TZ6Rog05+6wUdqvBGIUPK9Pr/5g4BXaPGxvHO63OgUfKydgj
ezKlHHjjsjLhToW69k0/q/NeNSOTvpTnScrq0m8XiMZ6nP+M69DJcZpU8OZCZzSW
RGl5TUCxx2Oemcgwd14NFBsDjPUVkGCbkCSazG8RBpFyuAOr9wE+wRo8qt6hAJOW
aNfNw4mI2OyRUc5Y4tMfRW1vAalfXfzW4LJ1AT/M0WlpFcWdlCTKEFSuexChNCJT
X4PR/fufdHc3LSJ5t13h7kYfZNrQJMr0YZtkMFcODigcB8ea0pbSbVz5XuF8SiSb
qq09xnGV95OIILyaQdzEukAw7oZmKs2b/sSrCYg/8yiVFc9tunqtbas/9QV4uQmV
JaQfyxvHlfSS1V9LajG96xZlMT2s54SARanff1vo2wJjuQFCrMb/1JwjHyYq1von
BH/bx5u6aDiOWQBT1fCb+SpcUDpkpubmjamMUkJlPm2OAPEU0oKmzsElvhI3F3Jq
oH9DK4IBJqYQG2USte8s/3jVg0PhkFL0NZ/zmDhkUxzvpCPl1eC7wb6pmVzjy9t9
RJYh0y9zCfJniiw7IL4owZaJzGVtVFY1WIfAATLHKcelMdiP3tQRB2OG1Jf7Zz7I
3wykhAWoIP06+cohyn76oiF8af1ZJbQdjYBzg9phDIePJcRw6jCOMyfGvXAa4RTk
MS/sssE9HBYc9Dl6ITTfn9MihO/k4qhSbfGHKDOqN3kFRBnNPkVfn7O98endLk7Q
PHM5RxCGvIBmHSGI0F1OW6HUsJTHOgR+peuE/EbHh6Cj1D/9DxjjqYG1DmsGYzvV
3BFYqenL83hQHmK/QGNWyBryme4wL8pU7AOdBCP6fRsIBTcFZ1CTR+s59ySN4+Re
Rq/RvwjQqfd0Wk8efSq5aLzYUiWYVet+avG3f/rMe2Bcg8wTQJMMGxMWVt43Ca4u
47FN370DqM2ilMtmSv7RAzjGo/VBNL/OWzIfaFRA3UD+E2AZjjT6Q6UeJz2R0jNV
rKQOyAxEEyg0iswmQLtLm5jxUDW8+tk8tJLlfHIo21J5D7hMDHLbrtEPCvM3HqhU
ruManIkxLySUK2jCIzBhD/fU6fsGa+y628HZnQtd9GB77iV6vrWIrINAJyvtoubB
iA71FfrzX8/uQBa2q9W9I0Mx5eScwxNfKK9hYT1Vyx9j5YpEei6x3xSl1aqPSbPT
XU9J4xwb1d+kuwcl0+nK99B1IX2kSS7qAqLhZ+a+1ctVjFJ6GPQvE9ks6+ytADdL
sFtvLRqTQqtanWgAZ+6+rZaw5THjGCDpo/bavc6Ytk/gZTr2zc0keiZrPTanLKCD
dBJv7cCdPOWqqbJ1iM/bwk4K3KMwRGTDw9U+xOkeyI/9B6HVhUbTg43UQVXE6/LX
/8PWAXNuf6d4vP6fXhl9+aBOJlLP/+Gdf+uNMWKsokI+wbkyG5OQQZ8BhbzAGsiE
y50w/M4A3U7UVLO9psM0oZttBDyMa6+HoKP34V1V8V0wBV1xo/s82pC2vKXmx18l
qkXNQsIT/0/4FN9eGPTxztzSso56RT1iAy84t20Ciwsx421CsXHIBQlU2DS6EWB1
M4OoPeQiF602a5WzTnVtrGqZuMQ3wv3xSsZvEOme4xF0kMOfzXHEsNxTWMo83S2F
lGdM8vW63zfkOz2qBt1w6fVHHf/SAKzrfEXlm7dA78T2pTIK5swan4+TsFJ3K1eR
skg4wusuSG7OGoCf3/7z0tQufjsd89lkw6M7ygrxkouKhUXopBNOHbNr8M3riBrM
GVTPbyapfV0ZRkD3toMYH6cAcDylQen+HPNdT2CiiUvkeRY98g2nKoInj/VqClCt
AxnozIBuBj/hM/MkEBUuSq/WjWwGT2HAxrlCMAv91jHTb1u+/ca4X+OLn2x3n7lf
jgoj4q8VPhwQsjn9Fag6CiKqb4i1y2+OPCfTixQVMtmPQM390FSrR+zVmpeCvIUI
0913r+4Ml2YHzj9u/6NZ6sw4SwisbrNWAxG3syiwHM6RR9UtINoQ/viaftjYP0So
ze0A0zhRfD+onk313jOck08VRe4viLsRXPtuq7b5Ax7HWYOu2U52s89aMMgi1mE6
GHxuU3OUQ6SZwcxTe/nWKBkwT4I0JPz15pQbF7qoCht1EFKx8AHhA3tUrt9nsAZW
1NlWJto2DEkySzKCeQXbqvZq1QCQzhWOGB8uUNaT1btAM4Qa6Oo6uuE36oZ1kOcB
qu6cF12h+9GFWH59AySaCxmIX7nNXydUOz4TjA+yPBaPacQp6ovyGtUofXouM0P2
2gFoqbIBEibKKN+iAwI8QHlv9bVyz+stqUgboGCJAytOZTrKmE+hEW11Zdw9+eKv
tzniWySIO2/EwiTjDlnVvC0yOckCI0nSmtQKQxAMKPoYqVNpC0TzbJO2Q7RhzJvC
s7fYPMgnt6cobWBz8PteG9D+XjkKN17fyFQVuw4BmzOpMglSJ0Zvr/DXeqZoIb6O
qq7cfpqldQotx01NPSsuUGcej4LQtoUVV8+dNlHDbJ9TxXkQYEjramranMfN8sxR
Hp0T1kHLTp9nKbCmhnYSXwd2VzsyTBDkWuH8dY6ugElHB1CXRDI6E5NTzdGf9a2b
BsJfC4hWz78x/RxqGAYVugMe92vTVAWHLkBOeXgFYbBldUmGB1JcJqtHpZZmg6xM
wPBU1wmvNRcPTcZtDA0YsnbzpVimmcNW5IrXpTX+GnJFbF/YG7aIcpGMxfKGzK9W
C73X09ANLpPWwMYPlv1y6/fb/o3cPiv4mh22rZdhEAz69xk3d//QiOL7nFTFQ0YH
Gz7JiMtWn3gaLkJD/3x8sfTsgn/nMo3JlI/njl9iH3gi0hluYCYwIBDJRjk6Mekz
Y7RLahYzfDDRFhYWO0VJx1S+yO0FX+hn66FbnQiiiQaoenmGYVwNqpS88szeT0jv
ElpoFjalkVqvRWt8pf8mKqCFXpCt11peXJCHq8PjjA3cYH/ylUtjATECEdTDFJrK
n8mER+72txO6GLmT+1JZF/w0nrWCucAyt5+NjTKxSJqZwRmAQbuvvXG762uEd2hG
78c+pwB31EBjggjOKBl8TIK9KAqDW3jgI0ZO4pv9m1Cckji7ClB+GKym4zSqWhs9
9DFNenIskb7g0sydahNBFud4MfLxjgrNLbhYBFpEZkHh58pvh1C3O9qEjJtED49l
ywkfhIL87zDqGQO3Nk70tNOf/dMqD1T0g7ZqwZdoMHs8UsTsi7F14OaAbPjG+Gan
97Xo0/RqqQsJHFxtSddFmkgM7HYYevt/sIM95tawxs8Rhj0/5/Zas0dNZdElPiX4
zuySiV2vi8dKAPc0eke9IExSGbCGXHD2cD9MD3RPs8x6us0sAmF8cNle7t7EMkr3
n+YPMNWtcXjucK9XAxaKbZ6ePb6QYGp4c5Y1p8G9ibq/dP9meZgegReckcNdLWQf
QOnosjzyEMCRlYgzXcSsOCPMOX7bMNjlZnTzkTUwdi46ED6VF4D7Y3jXzZDusD6X
zTIUJf0QtmhLqBEtmJO66FdcXxYoMlnAvjL1W7GRV+qTNPr3DVZZGsMLioNRlRaD
pvf492mf7K9XI6bmLL3IrsyVZc/gwuQ6mQSYfmpxx7OSRb/wzvZN3hZTlju/iSLp
T1KLq7kEhEJUD930/0T61PeX93stXdUgXAg1Nr+XnLLq+rtopkKF9MFlTAfkY71L
dneXV4UpJYw3qGt33akixGx8l8JxD2GgFkza+jNkv0S0GZkGwy6fEnKszV5Y4fOZ
CVD/gaxu2eRImkbxVBIqot4HN164zz+QhvLukBBgrRKhpLK3xU259KaYTlMJsZoY
Reb07fyxB2f4eNhr2B52DlXw3JuIHx9MxUI0W3bukssy+GsfMkVjeVxQzLiAeboV
wfgMBCEXO5zAAjkNY9UIaKgbzzdibb8kNtQcUxu+kOZ3SEqihl8aeHPa2L1jf6Bm
pRYF3Mk+q9Jar8ublUK+zfAu79SNkHsotyd/iLQSp16QamQXNriCjaeVXOm+m2+l
3E3k/0WXlklavlAj015BCX1gW3sEAoAnI+6zfV80y1kEuGg9hwtf0hkJhPZ0T7I4
JYm0EVVxB6Zh6eK/Ll21g7EuQbsv+TMsnpyA/Hq4XQ4W+OCPvdW477rV7MUpoch6
WGFg2Uu+lBmp7J4jASlad8htthsrygzPERV4SdxyAykS4sgMuvbcPZ7ereYaGGZk
IcPHHCpLoMogtnhsxZvDz6H2t+V/uRgUSbiy0uz3g2VhUli4Aqcnjqxhu6Lb4TmB
EN5KCHZuDv8+QSK67iOlU5EKHPgd8/NWg+Syf746gVkNYcDNXKox/OkVla+ZKcl6
t+Z3ONsl28UdijqWsG0QfMPAZJmikm0sv/DtbdHMfMKpni9Spci7DOGXKMu8Lt1F
WqOntiqVbvUdHsrxnIwbFdhOj0E+TF05T6SYj+TCxAnhartZkWRJ9a+vHQLkMYtI
bCAAJH9zOHh0s4fmOnNCdLhscz8l4BmbxxuzBxRrB8LTruNpOp1oguIQIXcSdhSV
T34gqXCtgH/GJnW/cZGGXZl/XhsGbeCh3gpuwI4oto8H4r5IyBU1Bc7vnG5wKCIE
+NAwt4M6gqID3He8CrgheZsxVQVqz+SzLCpIDhxcGH8I1ruQvCEaFXob877t0dWq
b5anIMr9ESKAgEJylIGSjsCXBeco5tdpm5n+zgV+OUHVy+d3xEUBP2ZcOxYzw6O0
m1FrLyt0Vo/AsMZxOQmqtkJE8kQjhSSOFT1r4d8uaCQPKhOZUPLSGvY+8cdwcIAK
XSvURhQyMi7ncAg1TVKt3JbEJXXVToNvptwuiSnnldV7gBkXxWxQmK2qfUNq+iWd
X0mMnYRPy1hcqXFnYrv6o8dXhhcHz4F9TuEjynak5ZI4owKxEwAv5YIw+8Vof+Ur
hD7hgH2ua/aMIX4gCSPqJspbMb1CkpujGCHErJ1ZxGj0QLV40VfP6f+NI/qZXy0S
sqiWUXgesYBk1Gq73rTAsMW/AlkyzoHQr/zTHsO99u3Ie8uAQvIXwIxRLEebSYPj
6m0JP3XQdoWyDvXfuo/uRPxzyBBVNxLzbyEWPRUo+NyzGZg5GVtvtIUnw4Tcaa6K
kOzKBSPSSvXOnyfJqfWGFvKUFMK5PmayP73j1YS+In73vPVxX0cBjwiKT89svZww
UCvSGtSo6Sj2PoOyQdhWpOsUrJuDfqPktsA7XlK8ogW/rquAIawkphYVTnAOvDnJ
GIJiJT4qWRLK/Cc3qOaWA+lIfDgO834kM+sB1jg790oK8P7dEt75wU+0ls/6/EdC
vYiueBA3NMvwBAgoqDz/ECJotEQfX/kfyVMuBrI8WrdjJ4Gi8M026EWxcBqtdNBf
lagJD+VEAmU/AwVJX0k43FfecDQ3NjlRKVScbcMSkv7UcpLpMgkv7t4Ueb7uk8ha
xQdUJNfTkLOwv48I271dsskNQ+QY62hp0MzGfAtsQeuCRp4oTVSIEeLq09LTz32v
2cEQObJSAjy2UdGXtuaUirK7poxNMyYlJQD4f9vjagYIVlMMzX/UmIy4Qy+NAlT5
xyHlp5fHQ+iYc9jyugn3g8FEAcXM+lSQyi7xJsc9j7NJk1XtXnHOd+c1GN3rC4u3
aV/5Vil8LUXtAH5qs06YAK3h+2nEQ8uRgwtOsuRCEHrBq2efNeshBkZZvCN1TIdi
5cSM+jBaFzFzdEp6Yvpi1f/KWizdKEts91mVoBsZ35wfzMzcbKknIbGWssHUS7+6
TBrMH6lHaTI5Ud2syCqOAPbenPzLRtewqePLtFkcwiNi1GHYrmOWafdK/U+IH/Ub
RHxkSQpiGfTVEe1ifKazlmN4O45nG/EMUJrVQznfB31Uk9zTyvj8hAiKIuGVyUVj
/mzVU8TCjGppglDLLEcz+y1dxpGlqdgtmXS+i/A4vbH8UhYfz4v78dfwnKyHmDq7
rG2If163uIPe5XYayBHrfnrBJQqxsdjopACwRHt+J72OJVu7v1Jy2TcLPOMZDl7Z
4Zk1fMuUqaeVJ3kdMMVT1IzGPNQPChOY/GCOKyDL0FaMHB3ed1smArRCy3GjM3YS
039GxwajE2Wfm6HPzHqmSI7ITe5lKJ8ZPfNn+nteMrV8usaOm2WVlnjUbPSipdqU
ySoYdhRpTcb8XSufIIFHUxmVXtIgoxIsf4DfF0ZA4rJ6iREfLKUjg4BCRD03b9En
uftiqaM6fuDAwdCnfFik0nxODuOBe2IWXt+emlLioWYBZBCkzjhQL5Aan0fdvS/c
cfnVMGiO++L6oXrjr5T8azp9a+sNEEhoCKKYcPqDBDP2nQO19aGuldtJRGFozVFw
UVhu2HrgGs6jNGryZ098VqCITmtIuTAReXNOlj0uciB4I1LUyjPvGvte6Zq/Zbso
OhfAFaa6RT+UazDlI6QX093YvQApYHOKTHrg+sbhJl3D/yibD7wwn6KC6n6P+gfD
/+KhWZI6PJ3gouq0nP32Z4R9kgm+o+vmHN5R1izX/34lML1+4wYOOcr04R9UY5Ki
qgMtW4iv5d1p7we4VjYQf8HMeCIzmc1lm2y//P/c5B9k6YVVDmC2FRPsghWsQfsh
sr7mL/LJ5p8C28t7Iez27h9783JtAYtm2Wu0gw5vk0fKdw0sVp5fnqTcGROU5f8D
nbPLYmTTb3jZXzod01h0rDZKbsHD/xRgxqsGTxzdUHkYNtPg4Thz3CLVY9TDaqh9
EhpbdXIaD8WZ2I832j0fCSoYeztfmcuF+ryvCPaI5Dt3hlYeBtQMwvDIBqr3jnAT
edl+ViP45VdjJDNVJLdRTyq/16oa1ALVN4EPtaSkk0bnNNKyOPs/REf3ukoMsTc0
wThJ2oodLXpkLPuXzz6wbz66GRVaUDZv1yDEgvyxjPt2aPhLXs3uXAa6mORf1kzz
MQdR7IwFZxv/fiY+YfLhQx/O+jqNmwxLLjOc3m5vguv06ngNfYUFUvoxwfJjmiHm
KzlYW6YO13vCVxRO0YvhBI+A94aPyz0ujqPxKvT7mCAkvfhluNm7MGLRyJxqSmPY
FAApGWEiZc2uZr+v+NDvv1xJqQwAaSd2WL4FofESc/TRQwizj/ihTMmZlWAMBnMu
+26syczsz/DxfK5qqtzTAegH+53ElaP6sd1o0ti0fQbV69F00YXj3a+W8yTZ83zE
HKTY8bVdi11JXsoo84O1a1Rh7xKg9QuZTxkOkuotd6QsFlj8ETGNGuOB7Afa7laN
Ghy+M8wrleFgS4tS7/UJdLVXtHY2tzW9TQ+Y5YWDq/tQsVa1G+MMSXC26v45S1vA
5SMjbSg5ychMvzTUeeExtFL72prq4wt80vpU1a1b4fbUb6rOqP9bv8xkG5CA85ol
R+ZqwZpXvfSWEROvEIBnMhKeqFQxz+3C4bdhNxqzODW95fKzWVhFkudqdHLx963r
+NDk6sEBYZB5mE3iFCEGpr5amsSPeaUnhtqL18TW0BQFqVySpuJC6QBs19FBEyNU
pXerwjZqZdZYPeAZsivqp0kJw9pRJ9vrQg7R02DeYlKxqOTyUq+vgWzIediPcmAe
blsdcecl96ylwzwiIEItaFlYouTGpkflPnoZOj4h+w9rvWb+da7Jd8sqsdFXfdem
E0rCIglA+sG9yPGPu8L0YKmAJtvf/pxBa/RO9vSvdKbz1nlqNHa5RQLsxS2Lzw6l
ELjC3aXZ0xmyUH85N6MGn7KW6luTIlP6KYi9sHP+kDL+8hEpV0F/OG672tJ2OOAG
CEzCvf7ocSIIEGMN4o2ysZJ5ilwriAGzW5h7ekeorvg5PwS09/KLvvn415H+09eR
9lAT+Ns9+lKUB1zJeTNQdBZORqSqB7Y4j4I2x8pi2Snc00j9bOKYlu9G7XdpEZhz
U0tFAHAaUG3eoKGk2OP5D70r0Pz7x7PoUO1LgewJ6/OHphG4fJ5pmc29UDWKnLQm
F6v2nYQDOEWhUDaqpUfcoz7Gv56W1zFL3W9Lp0DyKaSMv0d2Ee9zJZyf6tz1/mdX
SJX+/1yGSHIizFz6i9tf3jxpMEaxKZMWVOem/DkR/0g7W1K6VVL+Y9ozYisgzbYy
GKLE3ldox4b039s6WOtFVGUJOoyal5kjxfb8iwLPeMosKdu2xV/RvyAEb7LnsPPk
qm6CNh1W/okgICRtHcz3FfRPC7dOqjQi9dbkmV7m6qPiu232nKgX6dBD5wat6n9g
C9QI3IFUQnxgjj8fd+S9wP9jzqRyaRXeDM+I1aIw7j/7hEnVLXoIjRsmVlwASH7O
+Crl1dq1mMS0RnJ/EWQfQoPm9rhKhpzDG87/sEx/x/S9NqfCITYB0Ri9Ir4Oc5y0
ELSoGQDj2JmJ0rUiRMuf1+EVP+A/jZyMvrtZfAP3757/NpWR50QYIuqozhYGZDHE
M4TDbDYwO8TCGIDp9R3b/lDXf/HNBJKYbkmkKVNSRbljOlkQSd+KSzpFyQ/nB+la
K+GQ8c9aAv2Am5nhoifcc7Uv9K6sPy975SHYNfwtKNH9QL6Ig0u16tw6AqHvJrS7
EBHGw7cgvnLqwuZ5ZyJVBJZ+57p66T2Bdnz3GiZoojZMcunm3jnhQAhQFzLFETiV
o30j3WDAlCiVz6XiA9ijzVPSfi5gU8O1nkLp1uotqCkFAkZGXxeZ3/Vx5jXL80yc
UGF4DhnFXywUUtkYZIvSNvL6nRfomUrGPKF0GRl97Ky/xJXx1InhthPKVqR+7Q5/
DmfrnsYnj6mL1eCsbGUkpSIscm+TFDau+/DbF+ebtVxavAcxNWkfkelfINfnNYwU
c96eredUytX9gSC1/y7vdCrKJeoTEOnPN77nhPnj9VE0+SlA6XRkV98ox46x5UDE
27R3BPV3/Nh4g83VFT7DLjPqu/jFr61fPbAad8mc+5dcOUmeizpLbuXmJjWU3mgl
U9DE0o3WmyqUxidhHmzrSlUXXYOl/IMfaTG5I0cO+1g+soo8CIVJJJKRnhCZdZkA
NvIJznWmZ3otx8Sm7UUAF48u3XxTQBhbOJz7pHPsXCvjxM+5ZRE9wCi3R1F1BF2j
JMFxdTZANve0/sX7bfUtcEjdjEaRAOE/TNFD6lQwZ86dPP8a3HbYtVGA1RO42D9S
kKMIa8z5RCwPFYUug9WpUWkr3I/XrjvIJ/fW+N8wK+gSUfutq0U3O3Xo6vPLvzCW
kitWImEd1auA5DJVd1I92lc73+nz9S1ZTVH0e8Iqhidz7CruxOl/barpL/1dPpN2
DkHY2yOl3BA4os0IAKEOYOdIeJ3k3rwG+Tm033nhb1d8CDscdwsjrYOrpQVYX3kH
zYQ4WfQUIHMHN3R1TRDCeZyYphdD6M04ECSswHBkz3MtFdyoVDpVw7GkGkXcGGc0
E34UPof33zqyOZwxE1xvJx0tMdZE0hh8KGIVzMNZGYWreDudv8c1pG3xbb0ltcAk
R+FipKYKH7NDv2hgRc5dPRXSpNZXmc25e42wwdXRZs6+1Yxk9p6enPadmaWXievo
EZDM+SZCvSIy1NUmAFGA0OVgk5Y0vq5GAcslOdt8jnjaEF6hgEcmiHcXx+63bzqC
o8UhWNfQ7tiW0YtCfj7IBrSccUGlf01+bj+tnA4xo/nQWc5Exs++ikyQWHX172ez
zNFvkRYviwZFI+9JNou4r+l5Wgarbkc110z52cec1NTHlejbay322KmmSAOHcYGj
Dxtq9VrXxxwbUzAx584btJ82l6FEXv7sQV+VA8owmOOxAlNGqujOmmTYj4LzWAXy
J4vnv6n13k7D8/qgQWCiLtp7OLA6VzWL6xFONanfpCAKoTSdkek9LjQUkbA4gzw4
qkmVNacufxYgv3S+ZkbwwRvnNa/0758kMxOXJi75iGCSr25rtf8no/03hfAT6/DK
gdSBn9aq5JkG9d4BYL5R6ZKYdJ1JiLvA4QnXJMbVuw15eiSVkcizsgY8PeZCvjiv
Qb1hUpMo25rHCFxD56dw0bOUa0Yx0sYX+nyuA9CMH1BGugPPjBhcfL81ZQwCm39Q
McUSWi08g6JqkANisdV6DrDvMLej52R8RfopSJxmt+GgScj3Vua/HgcQrx95OQD7
MWlMCuNxU0Pv7+E/Jey5Qh+dZq2q8FyLM9VPST/BcSxMmRwRDut92pqi7VV+Bqjb
FyQupGU0GvfxPquXhw6wt2grLBAOutB/dcnszIoeDeaPK2WrbomN5P7JKapTl5Cz
ud3itFA1PXkmBI+JnEWImIyWpHEaO6A4cE2SrDh1halUwc9p7iEoaMEA/qC8votS
a8mUEMI9EEiDDtOei9/qMMIiZ3SKUCIdrE4SXDM09zZKL6Mpf32vzJB2JroDiIj7
pfxapymb3vNNXPp0pXaLx+gZL+vISXojMARimmmWPvOAg2f07aNkeNy0MOnnzfnr
79aRdElcKZ/sYYCTB54pqLqdvrb/tH5ywdVg3PrgvFbJmt9hTM9TlMHrDx9qvd2T
VohhzyyuAbxuEqljle3+nL7hul7DUet5oGsBMSOxr6ofSQjKvFHl22OmEdu6ezrs
ldKEjPfOtn6RXeJZhixwTV2zuBsyOytwBZaQ49d1aj0JSGpAM9hs7Uk4Tpzaqmz7
H1cbD54WzXbEt/r3O/qfP5nDvmMIYzKluPJJmNKCkdIKtLI7OWApsdn/eVzyV/nd
nGIs/dF75M8m/dBcysbX9I90OX/6cecQ69y1MrsJvahjIfT9w2zTSwKYvAn11EFS
XH1Vlw4z7Njmp85wvIjmP1BUG6BT7aa3OUkUzTqL8Lux/Va+rd76Z2lyS5SK1pvN
uDMKhT1y0rxQNJni7cyvKcHrgLKwa4pn9YpTW0XErw+sNKe8VELORCJe8x7OUzuT
y6AiBcJO9MC0xcCqnDHC38Nw7m3tQF/gcvDedIMEdg3ah10B6SywTm9gOrtsU0IR
+XEkbKjeg8NQpksPKAjpbnhT4ipEPcW1X6fOn6AkfpvLYMe87R7qJaBUHCPsuoKM
U2J28DiH4LiHP7PDeHiMBwIwySdlhYndRnSIw3uyqcr4VWBznYZkXZRrhBjemdzP
y6gxzNvfnWqJoITEaKYlZysdTnVuYGi9CyjIWqjvc5e3Uf/5lHPbCIOrqMvD2dhy
k8u9ul8hwZc9kjMjWBrWAXxftgC0Sm504F+4zsrxldEGNFhkY/wKifZEGw3fRFjg
dRUN3CnIZlbNZAm6saglGyklF7OHy5I+m6sqDkwhHbMLNXfSU/jlbD9rBY+JBrJd
/Mbo1ib82TI32+x7AgiCK3NA84o6BkRsMJ17tgChHB6DbFeFs1KzImOP2cs8O2Ze
jDDTDO0xSCmfmZpESHgL/UF4FLjATBysvZZpz/7bZSzDVrcSkc2q/7TC9S75YmDC
z0iE/k/ZipnxI1x8ZsD6NDvH52lt6gopgMnxD3FwciDNQko/bq2NL/8uIE1qwGNj
yES21j3IGDJ77L3KWOZbXY43J7+Ko6/qFFThmhjSQpKQkTIbMIqFUP4y/AfB8rUc
H6LW59ISjdMBawL9EZcMr591dSZH7jNeyi6rdOzejKMzl9QRDxtwm4d8PPb2cwOX
6yNUZjVVDbDy9bYo+qgbGgZFrPZLWpYhScNBZGyXJi0JGG132XH0s5tgHJ23ZKDd
Z3/FpqPLUfHP4zd2RG4bcDxWsUUORiukHxlQ9zV6JDxMA8OAmlu7MZCgyPVCfWtF
8U4jK0keUdqHrY3hcf2U0lVu27ish+4UD/bhhQ+AVjX5ZdPN22aFHnS0zTCefk8m
Z3BefnnBKPGrpDm9SVUbzWsSbabnwsvpu7j62Kmn1dlaWd7bbtrLRHL+3q3c5O9J
Ci91SQZ57lPVa887o/quD4gYq4efaLyka9DI6Z1I1RAdmfO4MDRlguSVNNpWPjhM
8IUWP5Dhd9pHpN9YPDzHK99Lj8FC4HKXMFd7hSHwq6PtnwihB7JvP6H+aJFnnIXH
dk+RTcqR1VXUmxG4w0vg2GXk4xwEpB0UOQGkD1YBzRKi7tZbga73CT/euzScEPbb
Uuhhwqvahv8GiW9gJKz/bdze1oLoxPk7ZPXPkGTB0j5ppd7GJBlOwTZwTIppy7MC
Oux0KIMsZHsYfsY9JO6WHN8hhXkZbyIzrxdopRijZ5DcUqs3PiS+wYjGg26AwKv3
zt39j0rdp5dOAyCsAED5sGTfY5TrWXFu7O/n3R6KcQ1nel7459bP8jJHcCG0/Ztz
a3S9un8g1JcP2w/adb26FQng2GcXhWdnsuumuVQs3XYrSNZxoEpG+yIZt8xdLdns
mbSmeRY4gZYV9LqLKT8Xema4FfPZlwjcHzvbkedRrj6SrjdV8zQ5dTGLzbD6wr2w
xgaSQervYWYtb/1VxOOEO7mPZmWpu69bU+OtuMmUHnZIl59AGIHehoL5GriaZVSm
Xd+XJ3g+NgUUk3Z0FnisL7dKIl1XtcyDAbUQgFV95VPOs8A/XrVth6pEaaFIPQKV
eoUQlHGByJZ2FNw9qDxGcNm4IfiAHeOw1SFGhHQyCtmc4K6/nL21AaD5XFq+KGa9
mU6xQl0b1K6HtmpYE+G7DH3MKWKTkIKX3TSuF8CQZGtEQPrBVTiS5ksioZkeDknt
aIqGIc5cTvxt0LtWXigxs5/cqTy1JNwPsiUPpYqq1xQe50I6CSS/mueDElKSoKX7
pjqJL6fMHH3a64OX1LANzx+8doC4r9XVieRQEhkXrMlwDhFYGPZUtU+oLE2Jotug
rPhvl4wfxx2KSRZjsfn/7L38iB5jzrl5ow/aViuIj7KAhx4g0SusA38tQfYBOGa4
URCbhN/D6aFbtHC36egMbXcJFzUu+1E1eTszwTOfcX/GkuBTfY0WfJnWgIo0tUKK
DM0P0lTk53Jjyus0DJA4R71z956qyaFgSccEeg6ng0MRTt6E0mG1Px8ukjEPQ8PU
w2Fb0EGvJcacilnAbkgkjKGWPKsDwKqgIVvjVygNiHCK3tn6T495j0V4baGBQPRY
+THsEn8toQ/p6AN9yMT+gUD+vHOP/jg+O68LQ1+HGXnAQm6BbBaim9yD9SuFOVH5
TfyK2ppRYDeL1rTQ+S9IpPAhluPS67eHCG2ka9IRz8BYdLsh92lWwW/OwZ0l7cd4
4lOZ34dJhYwqKzyPoxMVdbM+5qD3DljEdnk8cKZvaGxUG52d+atAeYgQbaWNcEJ2
Zd4+gma/k2ZRTkqGCuvyRudyeQ406/2hbDKYspFKB5b6bb6Mw5X06R23STQA9HkX
5bQ09wDztPF4U+Bj5aCaRJ4OEEnkdOr06qjnHh6qqOhLaPEPN7D0/n+xoPkf+qE/
JTfhIy9UDCb9SPfnpuOZbnSK7eaaKZkdY1WA95Hp4A7dOTwyVFmk3Gdr3cLJElk/
Uf0fo+viclI1Y3u77u4oJWWG6Owr6R0oLLBhJvsDuKWxsKvgpRcqm0apvYWGRUER
rGlfbjKQFRIPRFtnSJHHmIpgEHsvrmtcy3mtSYIm1eCwKw3ywDXtznfwBDv5IQcQ
6mT+wZAoClPPM7zan/ieu9RMaHfURBorg6WPKQI5rACpRJtRqTdyj5t5bgHy1Sq2
gCRs9BnhWa39sXMCiU6e1EhAWbEHQieo3u9WUo5U5iN8wsXfyJ2WkhpFHARVKTWu
enmEdOowKUo7R/FaAqgQB388ypjf2Rc0KgZUZ95DnEZrsx7p1PBCrVk7znXWFaUe
hBcYT7U326tzOlTTSgawOV/YMTIgxzLbPWHDj32LhSqYdnRMbMWHVXdg+XYP3b9Q
nsHv5oBsNvemJ6oyctmf4MvkPGxsaPG69K9utBd2E54YB4CAasui14nl10E1MvI9
8i3N/7zSLvS/8V0m1BHYJryXwqqEclN/9gOGQdm2usvJC2zO3XnxyksermbN8Wng
ni6dvbhtU+xFN/n4UUGAIbDBL8AV+IYm0LRqYIYNa2m6tbths90DuC3i+KYjlTA+
muiW0lbNoMsFtMInmSxMewcJWdxgW88K8bkMKTSwSHQPFE7Wed0HqdvuSDlPW+5Y
Ii807K+BrrQ5ti4x2IsgCjT770xF3swP2GIXhHgQt89FkHMh39gQUpPRLScA0xFC
GzABUOsGrB62VdgTfQs4t+tZnrqVS2hND6v2/IKnZ9DfM5k0yXTAdylZ4C67Pivf
k29cdtDGzE8mwMnLjfJc5r/N9Ec6NNwryIgaOmaid3tEMyo4Pzqqh3/Nfgyk2zLv
HG5NhEdfprnqB+aRYC3E/UsRtFEPOH9RojocWXalmhO5Q8otRv1OYukPkVE9iUSM
9Pib0N1ExgbM6AxuGw2faDEuwZVyTSIePKXD6nJF7lc0+gzkSfU5G+FQ+iwVXiHM
Z0+cxKSl+Y+DKxdmrFEA6hP3FZfhbB1G1ZkhQQtzoqD1Kur4LflnVEUOVmYMktbM
DEUGABIE6BttKPdN99SRAZWrXb5knsQzcsV7aKQaP5oA0hWlcz0DntRfakkGQY/j
lnMdxSlzTxOgUu69vWzTtmRmE0+k0zh5UvpK3nAMP3F5rBAqnwCoXgcTIUW8VNAo
m/Mn/tb3GaOUFCpuvSOwVnr+WQTxWAuLA18QOIh8R2s+bNsr3uYuj2YrpGOzlMyE
f5jC7vefy8a9WLEILCXSRTgLUtERBrOKSgLMx6UXhMuJxLFusGCW6bVTXtXzByoQ
HCFwVHKR2vhxVSff88wTTjCCtunTZji++bcaH8u4/f2GjZ8nSpG27+0ydheNOhZh
WIUKRwLli7FErdLLFVnXIae+p09ZzHSU//CQt1iwPX45RrRefudApTGEfrgR/wOq
rVv2gecOz/iuxSGxa0AINX726v65nLtHIt+MX6hUqavc6hmI59LSHwhAjjwKemT1
eWjZyGn+VxVSHWiFMly/pkP1A2NlKUdEld2hs0q4Bv79cMcNjxNPlRNLDTgkpsKS
yJVbqRunkcz/fjY4crktf/UXn+ddJHmKfGZU7lMvLXlxI4V3R2UyG4hfKbQqeJHB
9jR6uMg/l5eXJjqZmyUgSdouIs7k0lFPaaUtN3bZlwia8NhaIp9tJTnuO7/9sP3U
i3TzVHHTcbQCYNUgFmaveuCEMtQBXCfwv+y0UEh4fefmBv7jvdllX3At1t69GCqA
Q8GvmKMcKXZ3+cgG061iptayco3cHqublAdITOFspnU4U98b0wOdovB89+wZcKDf
ipG30HdMK5dLGMCr8BGVfR9paWux6OnZ9IeGb4ec7V+pNL2scGDuF8OiytRXu22u
8/QHbXrEssFnGLWzXRC/IZLPTc3MZQ5cAompxq4BGHukAbKpBER/R17TI+9bN74U
PldKORu7OP0ThzWykzlhmvcbTN6vHQ03CcbogTKObmGKsd7fmimkj6VbMUDZbd9w
UkMDIEoXUmPGWqjuvgj+49fC7oy/GR0HSnvrlEAKS7Iwn14y+wGWk/CCDK25p0ih
/W+uAfwmYjxKD4Bfc98jmLTing4pqPumDVW9ixEn+lZiBblX8Cb0FnE8iat8xncJ
ZYA9zmKzHdVLthqRhs6riLcq4OQdcBjDGo7EPyr4ekvdH4PRGEwPNfsI7KHzHAZo
EwBspzYAjMDaW7z2Fhya87WXWVb0OqRF22xHR+foyftkf7OMKhPPApZ9isl+jeda
ZHeHJ+ewdpY/3c/i0Dby0Ln9BrSji7g8YM9x9oBCDIZDsQRZpLTz5fcHkLVUObQ5
GG5pO3G4enB8gukfKpo/Hx905fVSUIVVQDdv6cdAvXtn33K48S+J0b4ydz75WLTG
czKlpBZmP/66seSjNn/mDwKTpgQ0wmDDWoftN0kozcBPRw+v8zLkbtgXOC9/wuKM
pXvEuG/FOdWf8ARPImZihtGVywY46FaPjaVBZ8NgiM2zuUUGQpHeJT4BTzfSFZu6
jku9vudHxAZ+8QPHVvkR5Cu0NIHQPeAjpzZYeyOjSy1vZa3auQBNTtH8mPLJ65ur
Q7swwP18dTZ+QFDBghq7wWQGW3acyp2hvra1WWLrx6XVIX6zk+vJ9BfJRVV625zz
/sbBadeA3/aDeG4ORpzlELrWR4pi95afcoNXXfMZegWMJnEcb8otkotTEnvdCfD4
JNoj6HuDaWhiigq5wzxtULII6+627GNEH8cSNXy/J/bdNxKTvZh8+go28VDowMb2
DF0CUchOhsTOgsKpgLetA62Guaptsq2qpTbeMkfVcl3glVhA3/7oX2X+ptdHxOCM
Bv7xojVr6ft+FMJPq3H3WB7xAq1QCQdEGDte2R4wxHbeaQR4qtlXbd/jBbzAtki5
YXAtD2ObA1l6lDjqfsW/nACUtOnWSm2mqE2TlxdX4BzYUfC0aKrJ0BgnM9F8MVzw
SulNJbsHiYl84v7SKj0J3ufe1+fAJRefNPp/FKQpeugMRFfsVjxuRWWIv8iDbUTM
egdHlN1ZFVIL4yHPNl2pDApR7yat0FkOftNTHtKv8J97jdthVaKIW9MEoUbLk7l9
4sHhcEI8OR84WL7SWBlbrkt3yZgIuymu8TCAplOevn/TlET+K87jNnuw4DKPYKsW
5cs5oeqXYqCPevuqgtkrqj9qRrib8M5ad7PJcrFhDEmna+PsBrMnc5tZ3S0rytqn
iGOaiuQjOO4yCfoP92+JTd2DwatraJ+YhIOIWJybJhqsFuQPw9HBGuqwszZdpo8r
NVrggbjhJSWo+LzqyMEGL8beF+PenxJdG4mhnvFQ9qJVQA5hzB/AvyXtvltw1a0V
NYmhEGrFfe0ncmSk5rIlikfm9XhoCIXifheuXWWmor2JEmTfPqmtN/JHQQqMjQ4o
EiBO/7oBbqBisufr3AEAtkNFMAIMM5+JjzaPUyaL9x8Lu4yO0ABO0LsxGD5uQ7mZ
z+M58B0VhQyVlJjgl/JH3sTPlmDY3prC6FK5hQsalRueLA9lnolLp5khOmmMC7Xv
C4Ooo6UdnhkPmxlQIDY/htnG6Fc65tU1J5wbn6YxroZKCcPNE+rUwpf4wlnhs8fB
+DN35QWCIzQSZ3pyAsBTn3Ctsz7ZhgYEBxWgoJyOJwXGv54DzKI5e3tD6pI7OK47
F9J39LYibONYpAQuiJASKdQU4DIsi2ckTpMpswXHQKKRvdfxSDACBaXYfBfXz0q5
NGdW5mKLLxEwBWGKyGvm0UUwEJl7/ynVCvEJwafa8t1mjgahnBJ/YIPsOkITUZJr
/OW2yhiVJ6S4l36LCTDwgFc6IFix/aSyabIEleLDZiadQC6Y3lGXlymsOSLA43sB
pctFTkI5gBIL62FG2dpSp+Pmf+TL4U3L+PLss8OniR+dJJCJLban4cBUbizcaXa+
MiBReBUzA3CVY0T/gvGnPODQ4MY7SeCJudLtFXT/LDJTIbE9aCnr2FtIVHPUkOif
4JQV6R/UJP/rea7z5w8cqAztyzptDLwejGvbf1p21rWfayfEflqexlejBNBOCVBN
4ibfjevfXRbsK3d2bXGG5UddZiEDaj4ANhN3M4Pw6KJAMeFPaOxz+a4s4r4tV0v0
NgXgG3mvlOKVHxFrgyfZdP6l7hgs+s1iLtpU76yxvGDPAFUbYaBIGeDoppNKWNCS
d9rah6xHfOZj+RfLbgWACQRX26Do3VhHEINNIHOskIxjdDPV/rBl+WgVmgXgvAWS
Fdlbsih/jomGpXIWTcRoVvZntLW1he8M1BBNEEsAbHFUKRDCX7m4tcbCICle3BYT
RRWIwYbE49zz5DQp/1msXznLcfhoXSMVzPUanzZWOMsKkjmzaPEUbgTjVwMFcgJ3
ymcQkr30X03vHwLvXC1HQwLYnJ/r7bPh4OCsIAiTu93I1EWOU2MDSQVL/gZnplaV
BktbOCurA1Snhd9Q6S1kVw4as+aljCNAInS9UtRNs7+eAnuE8p2ZVbp0vOKKrNId
hmYyqGhSs9tu4xVBfr1t7/qx2cQvttNY3qzc2/b6ZndoarxlAxlauO6eYMttivPP
r0gPJQUx0ygEqfKeBOlg/Q/bsK0HCfaG8Ny6Zb8uhSWg5kCIVvJi2puyxaOtl2s5
8XUnP14htA57K9YfYD0UpCsXo/q1jfHuhWQn+K4RR0SIoS/3uui6GuMAlW0GbX8o
cHqCTgdOSPVeLunA4nNqkjvlOYkqwDrCKizzM/MgrrXXYb5dUpFEr9DBQtvdhUzu
Kmrf/ocfpufm71lSOZoUs8g6rwTbh5swY9A+zhNl/NZG1XcqupZ/sTYo84B7xqO+
DiQd1AqqhjrvtjCULCzv+ZnlvbJ/QLtE2vP5IlnB7mYTDHbE0qxc7CwBbqSxj5jR
Gdj5yYOr6LfbfJcmxQueGek/ldLqjEVaQB1Lmlz0Jk9w+35VwN5r4XAAsW7jzs9M
kXbp2bnRTKvP5QjCtRocZAdavWiwn4Q3P7QGFRlhAhurfXhFsVRhvQuamw/8pLvA
Xrl7jOfRcBhgXOXdjdPw5Lap7/8WhVdx/pq593L7ybWUIhUIzOSZckL7U1LRzVRy
TO+UFypKbQQHasJP0oG6fSafUEOaNFfKFa/cE4+sphL3jtqVPRJ1HeGXKjvz65jC
cgjD+u6A40E8OMHca9fGVkqP/THXf5qwMQ4W+G7CTnAa5wVo9aM/QATdJ2G62+rw
myDKvHQ+T4weTYigSX3mVxk9CKnGK4qayIQg1WY7VLH540aYaCLfI1SaLlHsc6wX
GTeduzOs65j9+wQNa2aBSlH7ZLD9HdCpVqCD7Cldwi6abXC9jPcjtlT/qrkq9Y/t
I1upVdhkgN1L9AYfB15V39H207FkIbecDhS7puOW2867D/1+mZY0Zr2bszL5Q1w9
94EZXsRBAzgTWhpwRTfQ5lNMLrjJq9VMUkZVVZqIMlRAYUpul1QVZnGCaqey+QYH
SaQbTTcWZ938IzCjKJCEi+nBw4Tqj82nlRMGWIMaPqagdeOTYpC102A9cF2N3PvQ
qXnmBNUGdR94rWqcTk4kQ+IKV603LbXAYeOhc8cy+qD4qDoiYiKriBCGa8A617dD
h6EuhunLQU6V+XNLGB4l2oxmCwVRqbTKjwsisb6UfEe+g7veLrpoucz+NNqNyXTK
TPmQ8w8HkVQ3ntEwyporJLRp871QXV7f4/MYxsz8wtXbjQhXprbktU+CsFzFFE31
wmTrEMY7D6DkzdJsGJQXNvKQakIaljYvbHPwJzfpNfev4FB+8Chbj6DekA3MGtzV
PF2U2+re1OlIiYvJ517Q97KfB51bf25GIoZonHi3sCOVOJY96xSrHn1HoE3lI8Pj
tHcBm8InufZAIXNtHXhLUatxOfCIrbRy3muzotnjQaaBefOjhQM+tES6kzWbixsi
HoOgVkC16zPw2FwEajP+ZPvraJrbVlWWr8j6VGmokkRPkCaO6ScqhVOIzTCjuoku
iWOhGiELqDHpL6Xy7DPIK4RmG4nWURQXFHAktuOtihiNmJ9pxZhtCApDxddp0+0p
ErsEP6yn+5+H0qeDNbUrRBAB0l1M8nAxJbzCkHNHoRT+ZOdDH+OgoZjEbfB8iBzt
fOgVUewnJVojzovqcQavuxkAJG4JHmpbx+NoLfL8/5o6W5Mz4xfZ80zS0vciUG4m
Akx9dUMTWJY3JFf5kzDtH7YKKvKYlXOtKPWg/E21WwnqWSAdD0kxAc2UbWjQjtz6
GWTGn+MCD2nWJrpy3I3uAxeimuWMjG+zftNmmSaUwzxX5Do73bIQVO3cVnHSyC07
RDo4ohwA+ZY4PNT6D8Guh1tK5y2CnnlpHA745Z3Klq6lJ/VSsMcHaeKTGYa6b4gU
zbAkuC0P+Rf5LeD04z6yNaVArpzPX6WvKJ+DWl1YA+V3RoayO/lHkMXuntupR074
8WMmzPF+0fFDanTuY0/kjuMlXoLfk3psmAp3sUAJ9buQf0AeXH5HcvMmilkAuNHV
zYuTMpVVHRIPfkKD+5P/CkIlTksqlDX+x1cRly6EP+Hqufw8BxS9L9/z5NGZ4/HQ
lqhIhJ4Wr1fCaaSfg5aG+Br1Wk+T+2NIM7C9ptI0UE5lyDfUGDxfZK02MaUgx+c4
u6X2y2tLDUG9EnNp/YBeREmg92RskglIvixhL6zI9dYumhjrGBfPK6/1mvPZMlnK
uiH4y9IMCLktTZ5NYUmOo5MYccZ165pG70NY1d21brYqJBnFNCCbe23qS1AKUggO
fmuxV4+apSm/hVweivBslJmBxkBlgbRRYzZZGRY7C8Eyik8ZR7KJSWKTC/vQIZwX
D3h6IRp1/qSe16YvzAyI9wmM9joS2I5kxXJUApN5Ro1b7CbzIsXLlcTeTYnf6/OF
ZIlBwidmQTZIMCqWtVkcwV+Y6x08DGbHUKxQQuLh65bO/aNGdZo0EU+15z/4dERO
nOVo0/TgwSZpCuO6ifdtFx7a5upr7xnynQLHXpZqYgfVIPrfyFaJIq5+5B6Dm6wr
vKMPJGhNXzUCnVRIhanOMglriigJfHFXxswTf3d27QOYcVvZ0M2T1QSFGhgO4IfU
DLmhKrw5FByR69H5mLnjX2YFFMwoiG0/p88bS4EFTlcRq6/HXYtJZmNenI/IO+Z7
dVQ/ZBwnvA8W/FJzSu4KthKVPN+NhvvGxI50nT/xb2hRMcsRa6FASrr6iNnXvau7
AubVzzL9YgIJwBF53DqimuI0Zz2luJnUff8JlhmSy8Elej52lZHmwoNsS9O4QxnW
GNUFXDlkH3oXe9hTBibTDlRU35DDKUCxRrv3WI3TWYtDAhQJItCH0jUuyigzmScp
bm3SvP6VzUWkP9A4yvkR/8Z0i1IdCrfi17p57MF3d/eT+81OEMUmiRGAjTr0Yia/
OrXQ20WQPUH7O89QJgzPQa3PGfFuFyc72pkQUpQ+n3IIHIona1ZX+kJfUoJuXUCX
/dazKHleHMzpSKmVuR+RhjrOR4n6120IVSI6WM/k18Pp4p38yOvA0PYXrOrHLIp8
i+vMWTXF87SvhZecHn79so4AOxdfGD8Efhb6qQQmlFIFCWJ1jImfKqqnW4I6Iw+T
vVsGpTcuWGTtwhkBZpZli9IOi45tI+u6lohybp1DBwvEW6tSf2KrUdNWkY0cCZ/W
pxjfwuEyLQqmWL56Hs5fQ3wN7IKC1Le02JCAsAQE/bZnpF+vwdCl1tKYZtRGHW7z
LXeSqkLXEnB9iRwtiIkoQXs+pFpSP3loVHMLZdrFdEUIKLD1N0mAuEeWQ1w7npue
RFTY24lTgihyDtq20Ppp10PJe8G6y3HYkw5HPMgMSBDS2d5S4nBUmqk2TmMLMsGN
y8u0Mal0XAk2156w5qPCrBAO5xQzwmu5gAAcpBWpeD1niszrm4S0j9NSu65aurYp
/h/9otrXU84oK7qb00IDk6qWWHjeEpVMBRLQ0q9oDnUDtYTMC/EM/0OY9GlmpAJg
VVwnyGIauRcrU4qpa3hf7UO63dY6PITR4TMJNl93K03tKX0wNSwg4721midi3YaL
/YH65lJpbcbQekgS08cKIg5l3x4eSFTOGkbI7pCHloCzF7DCYR97suBHUdSYToQ3
pS3HKahnCRVYw/0GSlISP1NIUf923kupCB6xFIOwgqi66kKyL7kqbJ9AhfSioFmH
kyBXyq/ZUzKJlCqHUnpl+62UGVzsJhOEWPg39EFHECDbbU5kJ8soG1q0yDngpj4/
CaomHHfSTu1DkJ80rki/IYXcT9LJvznBSNEpnNbt0qR6bCO333CMOWmHm1jbHObK
YXXPYrpy+/3tbNQyrv91EecauJRPMFr+4CFW+Hp+gIPj/ZNcZfHcFeFuTkhoFqzQ
hKj5v9YGPewHNiS/fWVFWgcONgekEos2Lk3d7PfN1XCPVPGhsKJn5XETlhM+FF0L
ePiWBKYkqHytOB2gRBNb93J66H+DfLMbiGTviroCPILQDhRYW55OMnGrsO55PEYB
Eo0TwXBJR8PFUNIVSCM/ilRH535D4j8pESL/QMjAwmcuJM3GQdLXARHauY6OSTRa
dKR2rLvZjit4x+d2kgFaiaGlkFVxflDDLnSf7AeUKWf+zfmpe5cbPjBs1zcTrLQD
25YY49GTrxxDrCechcjU6tqVb3XGX5g8RZXTnNzWyj1SErswQN3rlH2RwsSlqnCK
SV9f9K31B4Y6WO09X8RLiMzSgv0rzgmsMQ3T+i4Mwl/5trs+cbQ0hvUc0mSQzA/s
8WbjO95c3NxhehjD5rem1rUH9U+9DMzIkLYZlFM2IR65f38cbNgKvadmGdXJLtC4
+ORC2vioQjLLaw8MpeCRlUyLuVqmsugswd84quyF13Jn/CDeFQIHD8xEi5O2Zpce
Az8t9NKGG3SrK0/tUQuGUb/NfiJiqQLi+AN4AoiWCMfY8KC4Aqz0tn5yrR2C+vwY
w85qzWS25vZ2gKYrGCyxX5LwJklTbPbS2G1KovwxR9bvhdkFfRookgpasGhCBFDJ
cH+SAGTetD7nM5TxL14Af533OcODup6/XLCQonLJDIh2rsqm2Osmaek968qAZrI7
A86JCVCstjuMwQegbcu1l8B1K/4LkmXhghcixExVDCei67u4ompdJiTg6pEyU4hm
2T+KGjrFB5yiQwCZMbiOtrOMWJtt6Rig5gCvgXseB3mZnCeGvyaPLiQap2AF6VxF
BZ4xCYhR+qIW51W85NHzqJnQ3ISZZq5BLVRY0f0TvazOb0irVCjA1LGk1kdHqEma
W+kfo3VF+jraDZ0XIZ1D8MtjenPJ7eoGhj+Mg/q2GPrWe8APGMzz7SXzLUYFq1pD
qDR+3rWzXvGU7LfY0+gU4z8rDCFz3MBfoR3nRtqnEoluBX7z9tnaRGuOqc8Fs2zd
IZMTlDbyQaIulfoyOMAOCNJupihZ2c9OnVYleQQQgPCW7lkDNnX5bXn8Ovyp2KSl
Gzy2Lpch+W+KkzleO7+XedRrsV/ypRDwtSJg6sBpVIGFA1rOy0G6eAssBxlFLio8
8pnOyA3FWBAPzwJgMlHoygKyeL79vt90r+aQOM7rbumUEza6epWmVct9WIolMYj9
E/kurRRLp1OB9b3X1HbY9gAu4RQG0lId1334oWdfDsmfD4NhMfaIWN0Th3s4nUSF
3Lou34BuZTJRqHbx1hUlSwNPUs7eIgYAUS6AYnA2RERKThpv8VD25qYiiWiZuaZg
mIkxomNusv0S8GV5KDcEX334s4vK+tcz6g8burCbi5BhQIwIcUzz4ltGfMmINez0
yBuyp23P/TT+rVecd3LQ7+8h8U6uqRP0p/7QhgGvnnNXSnHC7LOaSOI11VAuUi1f
v4ykfWXZ4WGYZwCzDDol/Jhrv8JUvqgXSGdLVej5fQB97ncolx3o3rwyApygws+w
VgAdtJN9ipmk7QKtA48IJVd1UEDy00iXYDZr+7LUVLmp8Chwfn9OwnxYx9JuLmSq
cwdEfHTY7M6KL8TQlBUMtyQHCSFxpjh0zTzH24xgKNBuvKfmPeME9jh82QwXxTBY
XaT7ektvJhsSuOcP4JKeOTFMJg7a527CXTwjDpWtWL7Uv0cuDihuQfMRf1nOAoJc
CEgB1NC05QiLIcb+cA6uFD6uNDOup7lGtwJvxqz8UvuFDbfI0SzUqCSwuLB2uCt+
IZO1FL+2Kx5AYSXmpGZ6EY6YtGny5hWWgmZlBsbvrQ6lYDqO5MtNv+j2UYLz+15i
Zi2CWsus+s+GRCeJfXForcWJM1HYqGYkCkYmdq4gEPw9VPiENygpU+ygmsOqAztQ
UNEn/l33Xs3YypW9c5Q5ndONp8WwkUa4V8BsF6I7ners3MPH9RJs41bUbPol4qSt
JxlxADUVTwur/eygmlQiH5kNn0gTvpg8b31QE0KJ0Izl+VArbWMBdG5tpGrkVRlY
wCqTg089CzLoIVBAtCwLhk98tjcz6lb4WTZkU0VzLmK0tNCJ9heFWYJig6Uvdb8H
ioDmXm/q+pzO41Lf/wUkeR1PNolPjgV868eYV35R/btjKnkCVcuU91k0TMJY+7DA
zPJBpt0a0xUU7flZLQ3Yq42I7vn/5El16ZZvq4zs8ViyxH/FnaJph9re7u4/tipH
Gq/tQWY9bz1lJHHAHwOlOe1KZX+49dQbg/mishmBhkexkiXhU13Fg84ne+SxzWs6
ZnMfhkGjoc5XlDIV7OjJXc6YjgCq3qRcZByayxM6TY1TjvhW0iOgsUUiFm7Cxw/v
dzesayOdGddB/1Br8WN7mbfFyCePwPUZu0yHtPtAPbVKTmdVd2DtLDrqQJtyJEiP
2yLu2oSFj6ZY+anfNUoXJfQ5+f4iu7fbzjZ5XV6N5YZEEwjVck9hXIkg6e6PUZDU
ccnCpAQllarldMkzPc06N+uwSSJsYzwR7ORZYC64ZPCuvn3rzebw/i7DTOh5c707
R2SIntmbSQ5r9YhD7dYIbGkUG+udO3Vfpv7yAVelOsvQUL8jcFRmrLhqt+xvcPOV
pDBrU9JdbPKYmISapqB36T3cVT3BAYlEglgOebaV8M15JC7BeqdVBhTkScY3iQ4W
kMksCnE1ZlxLZG7s6VjxRiFlCr0KZLiZLffW1sSTM6Lui+sILVIjx4cPEVEUvWri
lZiqEEje4ST3gpnWdsD9+fwDP4DA2z8yiv0ZFPLAOGkzfBluNPviPUPCpf4T/UwQ
zp2rnlQb3qaw9QUcTFBcIUDThVfRZ2O5zbo4bFok4LCwmwnqcMTeIZk1hjJPnfHC
lM5HCJDU6IZbM8Ka3pRDSmb1ddHDZ1YZQ0xAZ+x2TPM1cMLeNAKQzQbKVX4Vs6pa
uf+C/CkmFdohT+FBvhb4unJUxA78Cjz7DbKcoS0QI2fYIapb2+868CUaT9Oy9w/C
8CTjfC3CEzjwjVDTnqAgKJGUV8O7w2cDCCA5FS4IRy9Fx1BEmjjS6rmTApZEv4r/
KuEsRiTLQgJDyxh3Ion6D7n/J29d8UXDsF7CwcBSeIAtS/12ZoNbSYN5PlrzU+iT
PR1lu4wA0YSJ2946OOduDtUj6Cm+gW9651Pgr1SFk6z6OcmZPOH+CcoOW5nQG5J4
eUCD2CxVCpbjl7oLdsZOYAKQXLGcQi+uBS5odNJslkTxsoaucie3MmcayJDvjOOX
jmnwH8etq6MHyfrmcHLpKrn/jshPCcJWM8mcXte5AIBg+c7Uv69mW8CAqyGcg5CS
ZWzsbRWkpjT8BOwBv8yMQZ+Z4rXXmOHqoEQ9WDQW9jWMqOz5+AnSLsXZQf6+mQt4
W1bZs1LZTWWzwsSrathBq4R+T9GwaitcQIhMnvMDkZM3V6g4+ISpTWRZOB+8azBh
b5Lo8+wN879o8zfG554MeexcpNeXGQYaK5Z7dP37BTS58GkNUPpbk0Q5izqCQPVk
ohyhayvlHo4gritnsIdyouaZ5SOejTwatllW6gzW42XmypLv58VEU4yxcli4jIc3
zx+qjxsNBGDGWdqsQhx7SPCU53YeOXg6cxUGOcQXCTinT7OKe6p8LWLhIPk76oJq
RnshOHF0ksS6SHnhfwTYTF7/seAGa3xuBq8kBYb86T8dLzUvD68QQPdHG3j9jbMZ
RrGdjSvIjdSuYfn8yI+W1IfPTFsVFa8dWHjE4HJfNg0mz9FKT2A4DemS5R24ClKZ
XGo6aNFjzZKqEUzvO+oPnXEOF5rxf7BqQQ/O5f7664Ov8FVw7bu5vZk6QobrX3gI
OLJQ7xlBi7RFqiahMpV+/XjHBuE4OqS+aCpFnugEPFDPrem+WHbcur/3DvxslEAR
77vb/BckILtnOug2ZelweMB2wxu0HKNRy3A9glnNPbrryF0KFrLNSCYxW7SPgQws
AGpIXyDhoBUYfbE/ZYtNhGmgwyUboEuO7kOAH/VQlwpvp6YLfEvL4WOewdZqPaYl
1KXNhOpGvWScTk3GUtLo6t2aXBOeAsmlyMhc+pHsXN/Rz2I+9WhtaFthCO+nwPxR
KrTXv+l8nXlL9aIhrp9aHfQ1eO8omzz4jv8/5l9Eu6MoX6Vx3Zt6RjpMV9X8kWSG
45Ic1xAGQR8cHevAPz7VDCxoTuyPnCT+Ve/nwBohPamZ/TQ3EmkY1FHaZspb15mo
NENZKZCrDz2bBd11T8VgKO0tXj61lDDlrPdc4i9NHYq5qaUPwBgSAL9VwvhlXXOA
jaGbrK7tp488Ou6GcuyVtKqODcVhgDDTdcDujGrpzqIGSSwtvcboBDqvxmA87GWm
GMacn+XoIGNnvoxjLPktMeSwju34o/XFDaxz0iWUF5/unUrn8cZG6YAg5F1zYVeQ
sa/fdnARGRaIvl3uLdMveUq/qS3893Y6g6GQe5Hr7O4sEBzCZnfOsZSmRjWTQspj
+zgtvADP9aIml7VN3hw2c5Vvp8/b98JkR6l+9aZ7n+9/r1OVrPG5VjuaTAgWzLn+
CeHMZQ7eif4xGJF27rl8pYK8f0gTUR8xtL4gmisPxkvNlrN4AF5YOxBrCnabB9E6
nONsCtpjrdIlS7xmUdUXQc2V9tk3pPqlGHfI3kK/HcuKVd7gsqvEQCMEQFtpkx7M
8foMEgBaBw/F2iAg6fd1eKwtM4IaRWpsXG9jXQk9lcmQbNC5vfSjv6KUjHp9scrO
JSN4FG0O9iYqmgAKo83tqNZEcwhpvFlgPEoH4fUTuEQg+NRx+t27DC7YpCF/day8
12WdvcWAuWwDBfPbd0wbott02KPOoNcj4x3KfBkFOyzO/e7ZUtdVjF/RzJGVx4KN
+GZuJYwDJXdYhO+vwgsFrAWYZUmsLVq41+pVImqqLynBVzWeJzcTcOkcaZpYPjC3
+9t9hrr32iG7EPekj2jbr0z19hBAOq2Av6EqZfjpTFvfP1b9RFBzZIt0ZF7njMn9
/nbyHaoR6r2irXMLBRD4N5Lptk/3WMvhZ6gI7QslbF5YWxXbg27iRCZB8NoRuwvE
zdeCQlLHa5NAY5CmnioB2ozBhfDbJRVs1+m040ZguERm0RafebuCFejHhwtbYfvK
PcvFCSq4uI1qCwdIicagiMM1jHGmbsBwtpQGm7VaJ7AtlBqn2E6RcY+TLa0kYbLp
CvLsfNo4G/9xFmMfjhdCYAmz3tUcWWD7gq/FAkvSTAtJPwaRpMWDEUUrRa2Wmc9y
VRNoFy43l1uPkiGLwhKJ58cAahIXvRHF3Wcy5xacO6+Yc4IFIHB1fSPNWVKIzCPL
V6v1SuiBkct5sJRvEu/AiNyVypzGV42QbNjuw/TjNBx8OgMPOulAjj04suEjzVvJ
z3cbFnlPBnvT9WtoGiJ6FSxVQ0ikH885ZGUZXZBzkWmAuPwzspOI1ENQDOryU7jy
dxziJN7jjvX4UNSuBp1ohitKsRcm7xUMs5ZtIwqiRTGBYZ3JJyXcSKrpkWPDDZZj
trEjn0M/UkgO5bxRkmKOmBPbAM7iNqj7By9sVekB6fqmw//dMusPPJ2jm5+n+iHo
FBHFBsbT6l1r5B0GC0/+KQL9DF3Ug5EJXLIRkX7JTIW4Ia+PF1LILJxTRiVxGx31
2UF4VRWK1sUHxJfcNrHKEFQMji8oYZg3FZZXk6nxh6FNj16HixWt2/HsOQDc+IzL
OYwb2sI21kNRvInWq9uZMN77vaXP3OD4I2f8l3U9Xec9V9na8RAXmOi5Bfuplf8R
wPbnFWoMKSfTSVscE0n4zOPjjBTtQ7k093+bGZ4GZU2+Kiab2/zctH4L0p9ArAW+
lVBzpehlPAKSk/ik4103IWDGhGKTZm16IRrkcBsRIKfR7KQC9SBRrGUVMivU9OQ3
IJxfJMqi9ohrT6Mjl0JE6Ep+Ie1Kh4BDf71b1aODieestfWEtW6E0aquKSqqWlGS
rdCuYNUAJ+hxwlcDlc1d45WqCWQyvOTIBgcYN3HsIOZCTCjDz1U/Ir2zvTFNwdLN
ZWl2IhnpQG4VAH3sec0zR3lmIARLE92pIdQfhpdi/xrnEZo/7iYNkR0iBqiq3Omd
NbsEUF4b+aVZqZZX8alf1GjV/woqQEOb/kyc5bvYhcMTOB6wUEsngTv+fwiga3XK
RSY9RBR3QEIzW20uOfpGmZAJcMZVNoJW52479ZE6tZy10xRzkWCZx9PoDwNJ6Zti
SCyQTDyTLL1811w0LJ4Bj2ML8QNVhLJpnbBP3T8pMqeRj4Zch5a2Wi7S5zKhTFhl
8MFjU3jkB1DFS5M8ATIfiOCdIvw+5ByGj+LLA3FPBeVr4ydDNtUccPTv5xNE7WoD
LAotmbZLfE2af+juScEmV/59e4movMmqTY40zDzqK9ZOO2YgS0/YhsiyPjqy3ykV
AC0nSGtP/wNQWoPZUiOScQBlct4fJFX93glvnsCHeoP5b4fIIx1GdB6OMF1zNUiI
RvbJ2XOWMH9DuBx9dK2a77+1a0kg3b0bf//F7M9Q9CU6anBt5Dk/NnwS4AwSsO33
5FXDokC5/SMRsGj7Y+93V7S9CZGDjeQZVZCVIsB2kUWexqmMfDRykZaojTaV5BSf
6cd7p0gHOyvtDSPelPGiEFbfEcpPZozYdQm0dtgnb2gjKEA/FPbPIoRylGUFsatG
UCj8hS6kef8/n0OByn+s1p/bOGALgT4psxzRi8KHQMde6yS2oMKVzebE55sk2foi
PnZZs+t6SrVbwIIxCxrrZcc/XJ09GZOFYuvwQ47IX4VlwB2/WkUsOvd5akxRgmPi
evXgLZme84tMO5RZoqYb5KRz0xEtCVh5EXF9g0LRGGn5KtkMB21Lh6qIbJW8Es3a
IsqzDi0XCdSt8Mcr3sftfr11nmG8utqd/iqBMT/6GWDci267welQzJ+jQ+sfsuS1
Ubg0LHnNPgAaqcfJHmtycrg3DYbLAk10dxPpLcbPcu52gNXKVtXeLyWBscKho1Tb
9N2MSwUF0DJ9dbbkkfY3BzpR6FmpoA70tDhXsChcMTO+YtznFmXRpOQ+7BQiOjdv
bN5Im6iqPcsTHAkgggwhiaMsn69o8/GfVu83hbRHDIq2ECSKvf12pCigvKLFquoG
XSN1lL+bRuFKqALqqy1Ho0g495MF66UVg5ma4Y7tGJJuyaXQzQaMlAWknGIzCMIH
6y1VpyKqpKwqi94srZR5rlN+Uyv6a7o7xwfLd5H2nS/Qr8hkMU0mzevvogF6N3xw
6pj1Qfz91fSACUXM+qM2gVe0XySBiwNsaFrXfuE9pKHiZ8rInpzLN/huQ1kr5jg4
l/oNLRtcax7Oqc5QV/SRUGPdxZgfuruytP9cjxOhMGhPnjDVfZdsoRu3tvdisx1K
yInW4taL484ylLRiAZkqMj0CvvKP4sEhgSwI40dE98g9kQtI7/0mQcfOdR2GprBE
jRq28h1JHD6t6MoAfV0KICitcwEBFcBwkvhUh9nBoidrhWXLCYXE057CUrPaLGVs
IifH4UEQ2+kDsVW3d8tdv2tvpd8TO/QfiMRnLpadQwvFeTqC6VhbofamRoG4Hm4S
K74Y4P8aNkvrGRQgz1M+MqQ2WC86GrQXkG8Pg5VojAvID1TbxOKE3Msms0HL70Yu
SFgCTW1QaCm341783Yc69xmlLW4s4iwfbKytqVZOFuKcj9zHxQ7qVmtY+5174D49
OfPeuZVsG084Fzcbf4uT97m8HUIh/CsjJTOc6o5bz0MVAG1hHHntpjul6ExaPYs3
5SfTVGa1zAu6zhrcHQq3qmG6xMXm8oEQhTukSAePcEzz7FfGwEdcC+ieysoBqZ1X
Xoo73wGPXlZV4/Z49Igd6Spa9xvhPzIUAkI4+mymQJ6hJlkq1yDje/wkqEhYi6nB
bbJpzD5FGfpt02bNjT6s8sRim0EBYP0uWtBNyAjbdXe7LGJWDyaf4RkEkEyaH3M/
sq4yXlG5cMgBlgXYu4pgwJ/6gov4Abc/X+6B1W7sczN5GmDIu92cLnyXnWEY7Zxo
tK1xqze+g/IN1ZwZIzAtUxOXs9LTr8bBfz6OR7xvpY9X+MSZKBgwdZ+3/GoAMoc9
wZfOHbCnqWufOvckkHVoXIx5E/gcO+95FIybAuqEVdaHimf5TH9G7Q6LOcutw1K9
IVA/rZTmXBtPdvGhQPGYzhi254CW2cMvauIj2O0j9x9AgyDD2pwq5R8Du7ro5PQl
bdI+3+UrRfcALb438Efs+KNoLrg+6ECOful+len1ovFnRcvJQh44hI4+o3q0fzKf
148DjrRqyG9jb2i1qOUAZaHi7hzywQ3R2i/uStDmRlhaXk59AdvTlukQSYaTsBtn
g8Rv0WCFO9MyhJDuDhWtBLh5M/yO+kg+ni697G0gr6P+h3A2tELSviMb6yXrIrvq
wOENWEcozrjffL+tlvO9dA4PCl0LS7mp+RTMEi+OUH/V++FLqfUg+Y+3fGmfUELF
4PHKj47cMVSn7E0ol/4UB3mj01bQkvg3tr+t3wZJDwwz9K+fsCZ+U8qG7KjUIbOP
qw+F3FK1eeZjrac0Rkejki/0OJQchq2ZEyf/6SvHqHzQngzlgl74iN+Ermn/MSlR
wL9P8P5EjY4KDUWn11+/SoULXW1tbdOTTqvV5Z6UAUaFvhD0PF1xjV+O5thJeNjJ
MdV8lH3CcXJ8gqJYIUmaQXVFU7je3hS77bPwO8FvvRgQXjcMOBl/2L9HL5231CvN
dYlmxzSnn0p4M32c6uktahVXVX9STmwKFmwnowTQUoknvXid1pOcL2seSFVFvbG4
e77cIlCWbFuD5BgJwTAfu9tUDFHY3otJmyFjGzmB2wbTQbNb0bbHPk/CMNTL5AVW
YaZ4iNPLoEisHi7gGWoTh3PFbUAz4rg6GyPsXbtIl6UXF8hJjAZCVX6PVEoAJcgJ
6enEuwyEfbOtpxtpuW+cf34hhc8Y0gyFkRi+FEQ22cMVMUFpEKZxCMXSt2QOjD3T
GefZV0yB7Jm6jBm5KvTsG4oL/kA4DVxWl43G+onTkAEHeMKFj95evKEIPa9MTdnP
nxiprx8USclXRGYV6WBZ2NSjacJnDPmmLHUBoGC9LGr9qo7dGPtnbtInZXpeIx2J
omcvtYH2V50sZDMiy+4Qj6KdhBqy/NIiHjl6vLe1ygtfsflW42L2iyw17i6O+7CU
E+vMXGz8ySFQAu1/yritFvH/ERW0MhXZW6pJJHp7shlU8adm8ANzb0gGDge3qqlC
/BqbDQ3S6koyESqloRdBB/Z+iUfBxPAlVXcclGeRxYGE27GkQX5YSDQDCE8sZ390
xnaaIF9ZJZDYTqyKuwQK4edetrCSAjuc7ucIhePrD0TS0oxzScGpY7g0rhOPiYbz
AABOmZjpUXeorOsIjnW0ACp66omukJ7QUFTfAOagOQgAXZrIOo468x8WuItRLJBf
pkPyCzXO9NBNulXxnNVay+TG8beFjbNxDJvdlfXhHX2piGM4Z9z4zJk2/QCqaxqG
8wi9otXwy4uURtreqamCBcuLUEHBFMH9FY/fMHqXZCGYKghqZ3n3lB2IaOKI8pR3
w8Agnjv17uxH2qcU/K3f2B+SjDBV9GY1HwvT4f4lMCFFZK3FG/ikQnJEGC9cBFzZ
x2SLlYp+nRS/Xo9hMDgigOsx4Opjzpbqx4zLFas171iYxV7/vk71S5Qfy5pjYkzi
QMkGYmMrWux9G4woxUvCUNg4QISNozpiNS+89G2clGSHdoVQ1ERTQqnWcF2Ur/Nl
qizMmqU04QLCegNtCdEpkbghuYnVUJEE6hnMQRU9WPrZIN6LhOK3WzE6dMno/Gsz
mcbzhsCczwuN4AW9i8+TONDgrCTlHE9cqvacfL7pC29xs8HEAulBGYXwPNp/LvXZ
czwcI5UlzyvNqauDtUjFfP6wHnkTZkj/OwdogMQ05XIUZXkBQBFiL5TQ68HeR48n
kc3UMP/jLgNetnUsHOsf2UeMIHLDJ4Jb1QpyIdoH5i0KqltzLXTl450O6Y12CB5X
Y8rcZ0oTowpO9vXQ7RliKXS7UCYUJOUZz9yYqiM8xrUebmyFJjJqoxxmD2LuCsnT
O2pS7SW28JoGw3eS37eZ3Uq0BbEM5Pz2/n04JP54SFtd/Io2mr/o94gM+N7mh9Mi
xsTv/yiDW4Ay/LRjmt3udZ2WDfXEIis7nyGAzR/BmpBFyIAmdyqGeDQQbq1kUYh+
HPWsZ8UNJ0mC3FqBzYGPLTGBCHw7k3PE3UjuiOxc3soOTtxunCe7Ci5OAvYO8b31
nT+NFMGQHkXu+dIP9goLFf/ifCcXQDsiTX75K4dtrOsem9sAKHQlOEb7Fd7OXk57
5PTVqWJHqvH2JQUvEveKPCQgfjQWWNC5tz+UfmNgwvnAtorz9OKPbL/u1z1KMzP3
ZL5v6D4wzQbK2lfwdwe7rTZ1sUYuhQ6kvtkTCN7SEmkRnFOR9hnjQyaiT9Rxshjd
nOyFjlNd/uv7jklT6v4lYeybPgkx+Y6A/3fGadXV4Y4fP7haWbcjRMBt1yZxQzde
rjCe/RCkqEV8z1KNxc2gvENT7dFU+0+mM7plCvkoxlHbmDR0TQAqXYgPpweuBKMr
m1GkB9eowh+HjoZMQRnUTjGhpqTTqjjJjzpBun+RwyhcZipHfyvoIIpSeyAChR1v
u2kpitTBIOKI+SEUF3vu8QBDnXRWFA81ib6W7KBmVzHgg4UZlS2B3OqIkNfm4eSN
/Pb+rjIYd3DDHheYoQ8sjzHsBTckmI3oRffxzFicP5/l2+CNABljZGHxYiLbxWxX
k4gtsyaTRSFpDNvjEOjhpNTpnye1G8+JQNOqqz/ZzU1GyH4AU3RpN3ELqcz5GYOl
OaNh/TmmnR1jLrFHrccD7fMPqawH3PpgNcqgRRBr4NWJFCnqGqlSutVKWG4MW0lV
KSXEz6IVjSfCy2PoaBslwoL0/8bBo4CN+62R3QDD613/c0X3huGFxhmaJNZImfev
iEilcLXVPa14gTPWntqpp/9zgZR8FUyT7BGOMxtxr7+WibL5d4E6yz5SAQGZI11O
0uvw+aFm1CdUggEOkAIhe31mtEWloXB0MfukVDtm0pD1nqA6P6QAirtPamrPzKXR
PROpeH8n4Pz4Tj5G6JLB9nUqoaccm50tig2Wv2Hwo2vT8b6ds0Ec93RaDL11524o
PlPEVA7sAjv8p+0As3bJ8Zzn/hAkBJt9Yfqqu/YxolIQZuk8u6/SQvLLGvKHWhon
Di8w6gdRT6m1YTkJz66Gsw3DvnOkF4f5mgle5rHjm5eYJfxSSshLGb2bP/7qFJDR
UdCZoxt4M9rhuaIQbVaBvn95WhFjpK9ry+i4tBEBwpgTIuMNcwWej6Kf+fGWYqp1
qsOko5M7gpVDnWFESJcH4neHYBr/W4H0AljrFHJzuG70O/SYZSAUMGiPlXKh7fMr
zdB02izry/v1GzWHFcXEsTDaRA4GXZR4mgJzXY7duuFm6mKqRQD7XglgWD8fBSdl
FMp8GM7e6eEeqZfo1yRYJpC1hGoiAGDoGRf0fscVH9ijwjkivxQfkVFxI3FxLl44
wgBwZ2Qf8LrSLy+eG4aCVy8WjvXsbo9GOBD/254j3znMOMwdMkjPUAzaY4rY1FSP
uhIPXagFPV39NNUKWvDpmxYEPZlGGg0cjdJJ2kGbSfZZYBgsdLQ5tRRFIcs2Atau
tG9Wo7gHVn/rL9toi+/e5Hkg1KPinjfqi2AKvq7q9qZqHbLzsFaiGAEmBMZGYTmV
oHagMIkI+N2RBEv5cv40ajGvek3Cm1rTZmfdUw2Z2BjeySQofYtDPK7P9ANvT+Jl
ZNwvjwCCXgEjowb+Xylje61T217E6wDfPaXbX+MbAVmaxTWN9xoKKkhZWYr9SM0M
nN51KO/s67n9nLMHTwaWxjGHNN68b81j3CJ2OIXFWpUZkBQmcpfCs7M8DqS2jDTr
BPXx8DQOCf4HzrELTMWuoj3ivpiDUFWjNSAmbSOh6Zurj1M/HZtD+sBUKsB+cIeX
2i5Fc/2ZTNDkQf8w5QW0QMpsWk9s4AefXXVDkPlEj5iVSSooq3P2XkO/cxpy96hG
ZjynuJU8tb/eGAYqkkkUP3cGauydKp3tWF06x/CHh14ajmPgMc0DCog0eD5PmfJS
JY7/0Blt6zzH7aHxWLNXs05ynVXuEP8gGHiGUtunadrxM9r8ejuNBOPo1VrO/8q0
Cex8pR+2Feimk5GEX1tPHIACxHiYB52DOLU6i01O1nb+j9W/j+AOGBSLmvJJeEsO
XxzbK3LB0tEhcXb4GblOpb+2RHiVvhYj20vK+CqKPlraV1gXZmo4ij8S1F9uQH2A
RvCgsFu9j2vRwN8zDyVyv9RcW+dL3koYUAZH/hTA+LVgHmP6/CKM3DmMOaQAqM+3
f8xV/9whkm7ipK7zkfKgRVuRZLGChqoKd9MYyZJ7lQsfjYLo3yi4pWnhBfY0vWEc
LaBAJreOKX+EvZCqYs6WV3ur5rZ8oTAD/thxY9ohhCb+E/khGklwFaO0FjxmbxKY
Rv6G+VnpIvopA0QmQkhUrTBNxcXUjoHTxOy6+YrjP9Uix+ekZIiWRzoZfM2QJtC6
Nt9+VPGej2FEVCAFgmhHzA55GLpKUpX+/3gD56gvwu46oCPwW2hb5rUqOFlqxmgy
gZIiHxGlvw3kcUqYjTkPq6LKp39jOyGbVlMDT/PBBnx+U/it0nLGJ3Jq01ekTKJp
KxqCFgYOOo++1y1kDFzCE3GYy69w2mYAoGLosD/QHWw57eK5fXL4DSPBeWcR84bh
T1nCBXnNSpzbSfiFG52do+ZQthP+sHHRNsnjdqHXoFitxZ25YLgpdhVsPZMNE/30
iVfpKDnoeRdESmxrxvDAfrop3LMyH3sxixNceyeMjRBbp/EBifv9wQXZhKWL5wCW
YnA5qD4cLDHcWYn75NQuQazHd7CZnYwLU0yTURWGE3cP7tuIdIj5z5lBuKKMZN4r
FVOnPVOMxgm+z/LGHbXIPtt0jf5hyi3fjd2Sk74yD5PzsHOxkJU/k44+BCdUNWPj
SZ2ot4P+dnCS1+Xtuq5yZNxNMxeY2teDdbqZqamrZ3tzgkEyhPKmu47Zm/0QRv+r
ShpK+GHdUgYAXpSuX0njqPFc0xl4u8pdTBEL7yjcFSdxWbLpofipzrd5kmWscbYU
vk3xcYXnUmcjXU7w6HI9j1EvxZIamxsi/Xog+46fgBz9vHHgB3RquuvzfW7E6BGM
1KAuWfYsNVei756cvOmtPdy3kC2Z3cMOa6eBbYP+iTI2xdqN9PE7aNAeBT/5glPO
bTnG1BeKE+FRKFNBq9VvvR1g5CNvBuYYzPn+mg8N/M6yRxFA9ejEf6QXGVE/HY+v
+ybCq8/AgJdHNI0pxaQu3IsKFP2P97tTS6piW7mAhPPDoz0WoB76bKwj/ZywK5Yf
dYkm34tsWzJByMR8Jz6hqGSnMLBgbvxy1uu/O5rLSfFNlAuFPDbJ2yOegSSWDFpZ
hzzKphahujzWMNPMZJOkr8SveOB0ryLNn1GpDfLwIXTRjnzF+dbxpNOPodmBRQkL
J3vLbjDhwZFR4/f5BKGDqiX1v8TCyULu8R0DMsiU2YwcCKgFaUiIaLEBzgG7r4ex
X+RLE6JMW+mLSWx5hh6LHRBj79+Ttz4KN806bDPYHrqSqfSrQEbhRNWYcDkn9dZC
p7zmZuU/OmdY7qp70zAObcHs+udQ96oAmFzMPZW+xcIvkEPbFGqjdvxQKVDqLFZk
AIgI9FNACIvEL0m+3T+QauoWpZQDooD44IVqY8LMDOkhLsmNogNutxKRs5LzWkli
voNPbehc5+ZZhP6GuHFOzSm8rVLyAE0MKoTTNoJth9KXDxSBylK+P30l1BkBtptk
z/j4Xqlw5NDdcbz35G0IZWNR2ZnEObOikKyvJoLnVbk6cZCwPe00NbLhb6Qd8+9+
FmOTd67/tofy/e6rT9OIbARqNqyvdgA5OCLo4GGOgWXUBOzwnFwwnYTua2ejTz2t
yCtll0+Dgiazlwq80w4vOmSLL/TjfzyCeCqAlC18y5VWNmUZoK72P9P3VQ8QMqDW
2d7hoMFyBKJ0BqVQLn8SL3pM2ek2VFB5YE5cG/LauBCc8eBztqcdAe95IyiWXP5M
4NpzxDLVW10CpymW0oNcH0jNPOraaTBdOZgrmmOdZVB2ZNzgZBw4KXawIFUKYDSs
ZeytqIkntxOu5xG59Tzb+5t1n/OtBj08hWPF+PNJenC47Wg5ugMm9u2w0qydw6bD
uy+N+EUkzryhOL3F/Nk6c6z5B9LUXlLB8NSi7AaA8+NugZXMwaGcjMnYjjJyEqM3
zw7UttDOvS+/KZkPM18J3odRrG4xvPuBd60QTLHLXmci0lHVU5vjv+PAG64H6zv2
c41F+XizrWzP2hzMertlyNk85p0iamOOJ9oNADGFknsGXZ9LBVgPbyuR+WnFIu1I
bsMz5d3Aw66zea2JOIntv0vKYOmKIGTzg0zcgFifFqxDFdM/NQoWF/uirA51UEte
Mlw5CvDX9vuemBAcwJpVpp9C88vP8T75iezAE/gjrouot6+iOA+HAB6GXWcrT8hM
0eJPTTAyh7SWHopf+V9q0DVGvbpcURjXdYlPnFyVdPw/L7MJUjBR/ioZgh17nhac
cP62fLdOnWwPGfO85vVY04VDA0gadxtpDikA4Jol8dgJSwVqYm9ZjJ3YrWNDjoLd
PsI2Fo5Sfxx00ZZjJFTDpmDAxeSdlX43Colz/PVysXsMPVQnwnDOdnn8jZ3A/mOk
wqlG8KCO//iD8mKHhf0JaWffQKMEAG8BJX2EIQPqsj1C4pF1jDMUqb6yky2Cn4M3
IVm8Fk5gdPV3sePyQbpWSD4xrH63ziGNm4N2aBAMO2wWjbYHDIJ2mybIV4Lm/P0G
cojhP9ojgWVjXRvi9jANkEGyIpeV2qsVlY4N0vuwl3UI9Jfp2nM/8ZOcC+732eyn
T+Tb+mPRbWOCVBKIz8ollLvlDYItj/0luY/bhE89xfDpfyo9OdjKX07fpc/H7vls
cOa9dvlRurCkMH8MAOoJqCJNcDVzvDRiUMUsGXiH0LVyGesYe3t1wALwlFNF7NwP
UezfDmbpRNGxDyJhbD/1xhDx19eu1LgqWtVr1jRK1IYOcXJHO/oVDaGC3ODPmgXz
nuNt7mx0UVoDKHuY7urVgSCdg2AkIM0x6Ds+Ge/6rv9aiT1oGbWfZq4/ma3IoMoL
Bw+4UpVRUWLRPNhpZ+mU0SWRlRsYrWRx8oqvi0IKxEToeD2uwNCsKe7HZ5M59BoY
qAfuwW1P5y5MU45rvXGhnCKHG2YKVJ8m2FqJfqIWOAiC1RIyyWHt0pOkAkQh+bbE
tppHF4DXsdas055HdbJHtQQNYU6fHX38eICzPPJNabPm7/GPJq9vitK72OiI2DQ4
H0OzJ87i580Bb/Qkn2SaO5R7i0Mk1hjag7WeFNgi9CQUdTMEGHwb9qYngwMvLd8M
CEv5w2+nfsFksXkbTzg7/mI98F50xw2apu5nb4AfV4TgcVX56eegxSgJoScOQ5cM
xi6sfqdKu7gt3p8mdnX08XkF0y05bebHH+KbIvUVvbPTF1q7VJGyF+8k82qNhGDJ
sjcVmSshz5fXILf99MhPaCPqrxzuzoFds33qEDSRCsKH8wNbpXE+jJmh+niaa3FT
I+H69A9SwXsSr6eNuVmNQEICcq6C5XAHr62aXAg+ihNzpNx+7z1kEUizu2Yig24i
jQS9LIO6cXJ2o9PlJjTFGTBfdALQuo9cLAqnao6iRrfAwdfVhWt1o5ZqPPMHCvfq
DEhpdG0yZGIIbQNROCGUEyV0TVBES1Z4momGYX8GJ0q4Nr2O5FJfQQgrK2WecJfS
pfHmKRUe7m2LyX9HOKROT3T+saknrMVxGtu7gamWyzPSPoljgz2o6+TRc8xJfZdi
ww3kAFx6fauzkaZX6seRXuFBb2UdwqsaUTk2gBw+Gy3nNJ0W8s/WXoPT2hiE8boI
Yfv/gKSWit/wgJdgSqHd1a4valebYM1FjslHrOuUlNMnRg6wiH4aBuYzfCodKt5F
TvwpWpBYLBOlHpCGWF0iAaCakveEDVfnPdBNPesxH3s8p0DkpeVr3Vuqdpo/QMw0
0qXwJhGm7OlwdCo86VMCyBIaptAb+uY3M1umxg7LWQXw5cxGAGX07WRAcwOVF2qu
Kaifxdsh+u21kKnM/UtfhqkUDOS0oteXGpWZlsvc6ucDA3udUB2Q4t6CilxwdfTY
J7hc/bM1Bi3/6dhYw+k2uDeOxe6b1md3Zq+NYA3iNIO2R/SXYrPK5E25acYBJdoP
U+JDPweIjpwGUmtQBEtROld+0OnXrFl36fJvFC75mwGUJ52fAO3cIDhqOeG5KjjO
fo5F5nonv9aAjbaxQJvM9sEZQeorfEUSj5Q0Pxn7IRreNHZkR02GXLBAe2eXVxk3
52YnDipXLRZWCB6ZrdcKjAzhdBNSKyXwZjCH203QQ50USGomPd6SPLBnnTR8UxFT
AapgeG/Do+bHV809f5CO2AJ8GiyRyvxDVvzaeSWYpCgZDWW81UW4KigkLH8qpccb
9VHooyLktZRllvqBWs7MBHfcwJ+5izeLYk8pXd3KUlA1+W2yFvO3vq1hcnFKtgKJ
tD6WxOeoJKRU8igku7HOhlIeBQpbtgUn56fw1nmQd/eU3JcHObg3Nb6csKaKAw5t
9ORzL1HU8+mW7lKJEEmCICT0VsIFIAdAZGj+CNWZ/RpXR7RRPEsXI+jHVqTrJtk8
R3VNp3ZZJafyiUVQJi8XIXD+5aEemprndhCmrGs7iqLS0uLJH/t1x8xSObJuCMN5
ce1QtPw5QtMwOKCW5iNEGRx2BFbK6p3mKBonvoPXYplQEUAs34x9ppduDCjoe1FL
bGAkkMqx5P00C5CES/i+ysWBPkFG2+y89zhFJrZH1PivNFFhhYyzfK/RiZgnqm7U
NsosRAbB8Vq9PBzWm8Roe5t2YBBxbJR3oeUBjrNGFO7uOAhThNkYEiUCyDitz9dl
x9VXTIOcsEd+pWYMKV/afIogRD6QKSlc13NQim2A3A7tSOdX4mfEH9PNFfokfVPd
nJ7IJdD2VA4NcVyv4BxET0p8gpdqYlUeMiXrWcK431py1r/JURHMmvdIqAFRjEEJ
BVRlW6bMtVU3FWvisjTDS6ssyVsB97liz2aY85ltNsSp347GlQkO6fgGX7f5dYZn
8qqpGus5nblV2PXfsDqbf54veTse0cTd/9mRDDjXkdKlhcWTxUXDF+qc652JwMSu
UuVk/pb4MlvuGJEMHitXAI++Wh7fn4DPEJKKy1Unqp6BjW5KLypFmFXvmzvYNbcP
weZaLh6ye611YCqA/VTh55hkKKCIyBjotcDaVHrl3Bqvvdz1LltTQpIFMlVfIMd8
GJnuZ+VDbilMod5EN5tsud0YHBfljOOVdEDCVr1SIWakuL0VkN2YI6M8wBdTnxVH
5tVB+ufrHjxvGbP81FhnxbJe1VO021gvRfJvUYtJDB8NRoMBFULUF5j8Nujr+9VF
eQRbLc8JLDTljxLKV8OqjGJbS/0X271dYXYj/EHf7DjuxygT6QJYeSiGYRERJnVL
jyqPuWMxbUvkeWpg62eGOZIdeWGg3TzBaSbTkmVHNB9nycoVU1KBg5fIyEuceBV+
MzZcgIHuCiFmbl0TIe3RhAYOZ/inHDY6p+p0NsjVdssyr3IUFQeu33apLnSEebFX
MIX6sUcx1baAaJPP1yThYw4V/CWcs/fuAUY/5T3ugyv7dcHjcSra7X7J2OQjnUti
nld4mtRpLIGIqojQIvUxqa761nioJYPmMKOzJq7E9P0ii0TDrwiaFLxqoy/61NNv
BcwSfItBAaG7cHIvmvk+rS3hyFsO1OQb86dbMXxRoEsMnXfaeZzOsMks2zPJUHGE
JXS80cK9eH8Q3HSOTKnB547hbwPiljSKnT39rrUY4Ris1bqZWCDwZwY8hhYub5hM
LQCV9h9LhfnPiuBETHl/axYXn3HHzq2OsTWkGlBiYDMWPA8XU2l+JCpslaI/3ROz
CG/lTGz+/fZt8rnmAekD4MnAPxeDqEEbvofwHifVEu40Rtxl5v+YLn4qaS+fCroW
5HVcAxm6h+ix7GyesIR49Wjlmg1FJmxa2f1OF7Q/T35KsdODvb+Psf2EpO8cCrZ6
BTdQuJbp0ZtNKCZDzZkMZ6GPenaefWh0mmAWkUaX/glEQZyFL7FgtWfST0PsaWxg
bHPosOw1o87wilnz3G0UoENDQEyfbIrZzA0FJ7twvLYzCH/sq91SdKt3I97yEPpN
wX+mGnLNZ4UXF9sBjqo4heiWVaRz6ceAJjQ3Fzw1UCN0rPv8GlJn/b0ceUCf9EYH
20gpVSCfHeL2+9BveGaAGXwzsYZU4SDZq6Hw/uA7Ouqm+k3CLZfCBzkFTL0MY551
6zUW/dmI/J4p7siLFBJ4tw44yM1TxqnC2zfh7BDOj9xXt5cH2VZvKFCDR/ZBgYWo
IehZb8z4F5WXKQDaLD6mQyzOAe+zRTu4g3ab1Jaj8jAKrzsiR3n9hLE82BXbr8OB
unU9e30iP3ogoi8FUjo6v0ZVHBXC4sASyIrqpTWkFullnDIi4pRYhFXx+4OrQNQg
e55WizJ3Aihbi8dOYnVeiFc9YfgufeSiSsybZVnDPfQN+Njs0ibGECF3JtFCQBKz
Mo5/UbOfhxOW4CQracvPygUqgvjC8jAbWKBOCKBDD2IOPstiJXLgMwTpQnVt9nwO
uRHjFr1kTynmgy2CHbv0kqWgbzM5YkF4/Gn9/IX1SEpWedSxTLZitIrVEiknV7gH
gVxUJa28Y7/uqMfvY5d0kXiD84d9WjJ4BQuDFRn9es/LxeRBFzTE29VuuYYHnumm
ynZbGfgrf1M6EfLZRAXjkRKyBO3HIRiz1+WhFmt6Bd3WuAnAFVJKJsSzt6FVmdxf
LlrUAMynkH/e2CU4O4exyGevfkOdNqxaQK0f9raIJYCXWbqundIfMf3QS9qw8Heo
yQ3ytKgo8UWIZGmKZGR7tCdQER4EbOi3EyBgcquzeLkVLlOCC6fEAKDEvUnG0Xv9
HTCeAjUdW6QkLsu/CTONK3DsT3ie8y2Qpb7wndrWxvDc4/oEvjiqruh46OSjCnHq
+fWmElq5a+95i38+Sg2kea84mE6Eq8KBAMDd8NVEFemB8QPt+zovfYbSzUI38yOz
CI1Oz6fng3MxTSIkooJVzA6UgNRu/28WDMdZP4RGBTFdsPjkw5sG5lEbcH3ulAzo
svaG+IfJyG1EEDYT3i8xwifAYaHzvO/iYtTyPLq/jfE+0JO5bVD32b6mb3NDjHjH
LUiUept88v2SOa+JAQewtFy3gT/lPwcRK5czn3TzywkxqjMUhP7GAF/XMkXS3hTo
u3mWzGhauY9gd1zw/7Ki9fKsCWvoxxUChgICVfHUS2yNnVxYFNN70FwtiueuuLl7
pSmSlWQMnCrOIxgfYUkbGY6aRVeHVeL5N6BJdn6el41X1488MXk6X7hXVpOH00Lt
sjZc0ngDXI3/q1o21sYE/4aUrY7HnODTA/0LpA7A3ZlaYO7393YUGm+NEMLUwThf
SqsQeg0TKGhGQ3zNDIYy6ix0Hfqfcckt2NQoP62ZQJNQaGSYaPGg/Bpm5ibkH3bo
EqvMYSB0QQyJEiEfMqam3cJug++subgwbh15EZ5ScK636NuK1Hkk5/8rcv0o3aES
zuutG1xEHtTUR4poeKMd5+o6lW727R+J2BHJSZdlKEB59sbqoqg4o8jTxopEniRI
jJSglZD2WHMrJcbsPnr0TXv1m6EfmGXq7USrPuFPkrB+2pEptrO3bLQWnYSb7eJ3
OUincxls3afhDc2t+yj1lvHlWvQwYKSN2BxyWzdbT3Eit+TCJHfRSHKoOZwmG7Ko
VBmA7vW/7R7hffuv11DIMkj2XqeoQeaUc7Nv0LeFFWG6O9IiuDrcd7u3hTcQNRyt
R8LaBCodzEfocJg7d4Vfc27KmYkQwg3I5UuSVAuH7iK4/rxLU4L8WRtPmP7JADmQ
5KBVLiW3qdwDxr8hC/dj+CvNXmvRO2ubtfA93NeOb5t2u1tKSLKWelwJZ/G+cMi/
RcwJcHwhsicsEswtvnFbhWJxaTocmXLK+NZafpEqLOwq9QOK+Nla9LkD1vgu2f3l
6Nuzx5hTyPeaIUUYS/xVX1uKLIcdoGDQRPFd7M9AHXoy9k3FXQm23s11s8kfpmjP
g/X6yRZiIr9YDzJN0lK+pPg7oTwo7Jf/R9uOZrQ40szN5t1Y/+iKkwc1l6yt4WZq
Nvi6Wkc0fnZ2zNcS1kUw8HGJYdC/H0PzVNmE2dpy/ewxvzmoIiseXBGr92+mHn0S
hbiFzvWD9QAILyV9LMBGYSf4/ynfxCqOPHynaTaxgtZRa8j6EX4DC0aLGrPwHApe
/pZry4yqG3bguv+sl1nemv/6ouPlKl4HAdfiGK1ft+Bp1hcqsKaPAhpnt2teBYR4
h6iDlk/WFno3q9rgtWYi/sVzMKXBY0W0vaqbUOtaZNC83m45K30nudbVc1DxGO3x
dskpqGRA/9rVd1pEKD7zI+UoT0EEwQmmasLmFGrHgeF80tMXpL2heuxTwtggG8tr
DftrAOTHmuMb5K2TRyP0wK6pTkjPtqB0gpioE7bFCGuOoH+l02Bclyr9Chz/HFWz
YwFIshumP6jde9LYx1XpATw2Q5ozkPayrzVlcoAJNjW8V9Ky0phbtJ5gopYn+ni0
xwp1euqiFjmGnkbyALumxKCDO6WNLbMX2Hs5WUEfPt1UFXnng4HASUlrwDDEJBv9
osAAwl7frGpK0vZNfphUuvrBieyfsrOdDJ6rryKA4gOLBqRi1o8eRslpmyeoNCJy
NrtvkF7JektMy7Nywng04+I3N3KwtnRRxn58I7Y0wHku2sVuOJuE/Vpit3pAsS+O
VA/fOcwKYk4OgEwRLG7si99zSj0SY/qjhzzPLXYKl32lUUrHQCvxpLboZrOE7+sX
DLdlgVQpujYfuOSn3uuZeC6MOzkmic5uIyD/w3A+YnYKWLi9UzzjAGbzYQrQhPLl
H0ZxisPfFx92MbWwga3XtHBZTB/EYA9VkqHs4gBooQZ9N5RypZ/wAAGJiDWnmebA
TQBlRKNxVs9LOx/UQr/B6bGppDeVhZLXGWgjufYu1sVX7xOi3FcbNXIwiosu7Hlq
iibK3YR0j9Y2cl+XHEiU/sGwTVQKKsJBdc0PP7Bfow1IuBMKnSgVtjouLvwVzUtN
CIRgqKbwSIWo7M2UdOsAVzaeN6IU2qRXSV6xnL+GW7l99cg6SvHyQIKU2QqlpIUk
g6Tv6qEaSezKA1wT8lVFWMcNqV43o1mWLqglMgjtcsTVzwU77Lnd246qrz6Rv7EO
xYdOvjIAtI9dXZ05B0LUtdxsRmNy0YYTUJCOdsQ4V0n3sE66PMicBFhsbqN38oWd
DLSuLLb5j6NpsSms6ZOwyfb6bCwfUfPmhgo6jOP43GF+bXGKq5YPHiyEIAwmSXrc
IMlZfBkeH5fK3MNfRxniyrdo2SOfqg0YjOL25X8sXSEcAHTsj30U/69knqOGUuRA
oFMwmsvY5cHWQKWD5lMSIjwe8ygKVqk3pgZDPOLYUCM74C53YHht8iAOGd1qwbvk
Q7YMImkXtn8CBn+vwNp58r5/oW5dxpf9vXl6BhHp6hA3dytx7K90LpiVqf7oYwVn
qc6LAnOMUY+pK03Wq01zTRVmXiOnioaB4QRNYa1S5wLEdnElMxXIkfj1USnebkJb
X206ED3aq3898wCHtyXT1TIjR19EMqNSVlrpwQhL898IvxnCKe3JNlEwZltoqZ1d
KlKUveveuq9f7uPcDaZJmaBYh9bDabYC7I1l2dB2YwreeXx97Zhgf/3EedDELz+g
h+ffJGvQFRoebl11Kmsvpcw5QEv6B5IA4WVd2MD+dQJp1DYa/PqQA0XEqEI/yocf
bhbZyM9xognsLJQCXUKQlbbsbHDodtJnGeoIIywzQA7nTegl5KBWB+ALFWVBQb5n
0WBCLyWItgwATG8OJiAfRLdITiXwIyBH+EP97J3wm3MvpxWy/MO3DEmxWziECGGC
xtTIqv6dU8PyMA0H8FfARIwmCn6LrMYWJ2KOuE0gjXGoAikq2F3Ky/QCA1bWXL+Z
E2zVPX8WpqGqb0NYsUSQCmshpvs77LRjJuMTgGZGVQqqdGIsBFTM/XJaVUu7STtK
FFbarfpuXthkwgRL68AGAoj1RinyEd+nDLn3ldxvKYi9zi2/q7QMaDICPAWxwVbW
2albGu2Z7dNgO7bezKaBRmJwhVun0P+VbWbhuPaqCLFI2sukfEYhN/yaXdelXDvd
2tAc3jht+J3B9uSB6cVeANqM8ln5dki9Cc/H7HcdumxEV0FBpyjf6u8NgdZJC72t
ASLlodEUVFs+QAwNWMedfS7adU4GE+YH+5w6RG4NrHPYBDwuTDs4b579WL+R4Zly
Qvx3e/oF5WDIKVALImPYiXu1jlyt+27OJ+rWiQjcrFnNNxHbIQ/UoBZpGaP/bGj3
npSVFwLVSk2HEz0o56mGZuZKEIIJPgOab5muNq6E/uqiLU4HlzFnPmTqeWa44XNq
uB9MPHdA6R/nCMfBeY9c9AVlRhdGoI4+pb7Wk1afNbTG7w2ON+GcHnmeABC375QM
1fimVSmY7qwzKgocwXwXlen+GQCe8DMlCHh0yjVPSVGpM13p5XDmt+A8bXifTtW8
vy/G0Ub78dQHthuJpfo9xGNsxirzidFW9Vkt7fMSvhebVFm4pFGxbTBCLZnFKwLT
Cf7ZTJeskOYZ+bZeU7SaIuGVaNOX41RhU3bB1Aay3XGqPr57AbQiXr1OCYoufoOm
+8yMihqz1He7AqAvGf5fCZ2rGPZubjRfqMztfTMJOxE3u1abpSHIgXECQaLPA3OY
/JVPuHC3Zooo/ZK1kKs419ZOTMAdEtwNkJwkOpcrpcNATMkfuX4IvE3DaafUbiUH
gdtT1/gzuOlrNBh8RVMf9CsBJ+gRtcp60ph4EhbCM5vZ68S5cMFtrgl7v3pQgOUs
e3INUfoZiiGtoUkehpe6d0484ycLx9PkD7iIlwY2dHQaRcdGzTlZv06nspjc+FBT
rDzJPrTUDQK1nQDpLA1N6n99TGCjTbHLnSuPX2FZRP2rg+sa7IPuxFY/Qc/7+K7/
e/c8jcpDdGduDw/O9zosgVbHaDhLyB2DiLul2AGVoXA4+acDqHdm+NWA3Z+jR4Ic
vZoPPRFiXvKdlDhJ0pbp9t3ail296H1yrvyCMIR2RhwfeHHzIIxVSaz0dJuzsEor
rRcXbfK7hivxG+Zx0/+EMdvtEl3+BJrsJMJNx7TpbqXnXajvRnIQO0+gtuFCJg9v
Eag8xEfpcE9A7BwAVZ74oUWRi3MTGaBCsw0I6Dc9d0uNghMPxueRsbUljs3FDyPc
elov4XoEsaYmFUxTk8vctE9oLaGDrOC3ZkxxTWVQ1H/MlBrVMZ8gEVqrNxThAeAa
hJB6n7UkZd+UZf3fc5ynyY+IAWNKn9vUtY8Q/hKt1AUWOTSHyY3Uh+k/vAI53oFW
Rf+zbe2kVsXH2vvvq8JgiY0phdY1tdeahpZ//f8eTs5uf45OG45jwuKsH3PajLir
KS9UoSE0esENLN5/qLLtDFLXauI0GNKOXnujB7N/PM6YVC228PDZbCYhOfplZJgY
/z0g1DnHgyXosnDEZ6YWog2edI+R0QPPaxaCGeltIyAp4qVSJaxdiZMH4BJQRNhO
ZrbxAlyXT1iCEbC3EYuc4GD0yixu3iiujPMdMXSbwIDRU5Px1aN3+u+If8igvvIr
ej29EIFVGD2a4UbxmjiLma8TrYoRrLOoPk6tlXgoqGt5nIB7bpFS6l8R/bFKwGUF
Y8h3749YkQ/Rery24cjhgvQnu+NyhMWotZsZUoPSxuaSNqM681s/279EFxWHy2+u
kU7Hdco7BoQDnlpA/ztwEh/K6zsqAdl4W9zYBh7pvizsSWzlDwe5LZ8U6G9Qqs60
5cWmERR7lRtHqAJLT9iJ2WQYwcoES2w8K9PscFrh9ph2oOJ4J6dDXsjx9Oy5yhfA
V8s9nPd2evUta8u9z7usF0c2bFYzwC7t/iShkcPF0JM+GVn6TIKhk1vWQoNlAApW
6u8FzbpD9l+p7fw5jk4DiatS+NUUtrkdgPgYgAqcp+hVBIGIPFSAfhnKVH0W7td6
/wgbcbSHRKSKDxjHY4z/SXoj+biYuSEZ0icJ/HTgUrk6h4gOwZTNIeOEgigGe7RD
IO0nGkgdwRRPUgCz7B0AKxd3QvynfEpUxA2IQvVcThGFAE9qjPzeWuPqiEhIo3PY
cgdu6iOfBrHHY/Q+eq5eWRbg6S8oxNpjmNSyCSW31+xhvSlv1fWjsQ7jlPiURqDG
Yfok82yaayPuGcK2gPaTAqlJ6O4a8t0W++agN42wNioJ/3/xdiSuFL9cZc9yvjxz
u17VkHlaNlocvYRvlAMgonh8R1/QnBv3wDEz3sfpa8eEc0oPsLevFwSad3ykTnV0
jH8h9BvO3IKHkJvSqq4XxWiLYo/jCXEo28wnhzExf6JbmjlrC35n1hGZhrL3pGs8
NLhMG+cKcu8y8t8iBqkHMPG/GzUijy4wdPSpBPGmFejEJxVtvB3PStMjFPSVBkOk
OQOPFFfBtHUZvtUH5emNe3Ml6erB/1+mPmpfSXjdbALU0r3+725uZt6MRDvFixmu
fKJW8P2kRlEMuDg5Zpj1JDct3vpHQ0hqTcI99tAbH6qgjtz+cRWLA1irxstvz5d9
a5w2Nk21vGAa8sXjdUnvKkpcc9mSXeKt7Q1iV6s7vwU3Jv9WzR3MJtTPfi79OumL
saidTEzek3At377SUcRZ6BFH6wTWJa+yYtPdAZsC2futA7A4bFVTZzYVC6r4y1IJ
YRTCKUkVCB9Mhjn/me/ve+UZxpK00ePi5TjTywfHYhqPAsC33TWn9D6KNb0cafOk
sHmF1hNq6OdwzaEvRzQqvcySgvchyxURi1eubEl/btztrAJ42ucP7+siLQ3N0q4t
2kAiVqJlok8/+rdt6rYZm5d0CWaSyqktwy2LUSNvogi+XHtF7HJ5PjdggF1BkXHk
nBVNvOhfCaffyDEpOMFUpvtKBjRQ28uXuCAjltvW2pGI8BGXQxC6b/X8BdflB2Ac
WTun8lCf7I1v4k/TK+z3VqLfAAgeUlNIqDLJc7w/UIBfqdEchDl4FyEj1Wk2FKNI
n+6u4nbqVh6CtOF1AK28aB+hIghWP7JByDXD6o2r/kPTLqOlTXz9WwZsHr9o38Ju
6481OkN6TxU/v9ois2s4OG/DuO4levZI9axUZob04haxyYATht9u56dtC3e04+06
ut2nRED6O2SxGqXNW+drdTv4rwGFevAsZfBcU//ANq4p5GyjiyqzmT3Oqb/oF+xC
+DC+lJcUtK09NYIeKTKpti9HbPM8ilD3ebwr9FAwlRhf00bgnooqk3RVUlTcShi5
ycw8/QSKAaLwyxgMybKwCTAjyLNnXEN42+c1oGK5jcXD4u1sHj69+X5kl3Sljtlq
Fq+QUyA6vvAL6rn2qghIfp68e8Lj8AJ8xxQkbfg4NelS5cMj5ROBUSXnc2LqHrdX
PtdXVEMm6cV72mVIUUD3qi00nncc/C22yWRPFP+wJWXWOJflS2uF+ynyquSihn+I
7Com8it7Req0UkQz9Vz1nUAgkjEJNZCyhoae5JGv6tC0CmNuFeehjXqVug5BiQu8
3+nwlDWia2+BvUXFzS+PXcBaKJf2wKU6fNLth8cJItawJkzjzswyzal/3EZEF+o/
/oPdkyjEMIMGe08083mLznhfwUNs9I1HnBYJTAuxCoSpDeQixCWzNIeww1Wwf0oL
7b1khtzI4rGb4LM7us+aSAESACVIMSZgNyIAWpcVmLhwpGpXttn2Xd0U1tnZsNVj
oeK74SFyKuCfRnbr/ItlHG5lN/dRAqKbSEJuOdsA9F62fFC9D5Bkf0r64XVi/X7g
NyEj2yZR26suXc5WJOLRNizF993N+HSN4dc/9AivO13xixCmu8WkuJ3Gmlkia5oe
ij2AWl4vb4F7SdvdZMwdzyqvNJin2fucH1bNDrIhCKq8oufF4lFNVIx3OuHf2sl5
5w9cDxZyeWFM2FpNbT+Jmot5hJrXg3T+C0Ftv8tcHPxWd0K2YwIMGmUShmK9Qntn
MOYi8miGahUuTTw7brq63zWSOngqnq5db9+JxCwK4vbV6zkGGYiCSTbctVGTcGsi
JKuIiWDTvd0TGKwq3NuUn8NJOmFgqgdD+w4nUkmgOCRv3Uv/qb/97zEZyhsLQbi1
+f/fayFa/WZZCfA0Gan4N/O3sxLoJe77EmYk3EX8sgxG1LAPXKD/dQI2pGZ+Tkg8
jyxgUZHoi6pU4WhGe9+Asav91cDA6c3d5W7EyK8H+B8acU1pCdYq4fmg7PXnPu16
1hiSyRQbDMClEsjhwXYWTZHwuHnohvl3RfFWQ4mJkwtwSE7WI8e0mOHTZdqQtYUU
GHiArxgzGWRCT6ZSeFDb4wE8ppemiAFGpVwfBP6JXOdROJEW82i95aPNjoJEKijG
25yoT+ys1438XXnz5dlSbsIaJJOlwccICbIuMWh3kOaJO9Vkbp5qV48gEK3QTagO
FUkpOTA8WJRsotvtgFmcJjSLclWlvJc/OUSNvmgntPCQsp9Tf40PrJVludSa2xYx
/yY3QYtHYP5xLae/Swes/pwN9c8PabTbmibKdjYZvfk4lbm7ArlGhHbIGtPqwYEK
5T6aV32eaDu7g6R6sdOKyMd6Gm40E+v9SkakW4e0QiRm9wb1DLdpEdIYVFQLXItt
RRzI6EzPZdIoI1FWs7TOCHwt3ZOXq+fN2jGt5Lf3xGofigKHTQvlObk71dyp99I3
FjuOM1EAoUb2IY5aexc+x3yEzd/Ctkg7uyf1HTHYG6Cqj0FcfY+iAu4bsyfATFp+
RZ1A7qkaEhE+/92bfchZc7KKFUGz+IrrgIR3G1acUNkxXqW4Lyx0CER4/fLV0v/J
24XebAhl3QMB0s9O9517E4hU8gP435MQVHpIS23jPyhuUAmYn8YQcnIXfGa9Hr5F
Pp6+8sFhInl59Awwilx0rX28Dh4i15B9KlhG9kWmOMar8QnCBK2sGr7gD/Ci8vXY
Rj/CApREWSn9/hZ/eZLz6psnEbtsgYH3W0kTYNR/cUAp/URm82cKKQJtgZ4U7q1o
PhD84WTr45IVwoqOWCGVaW7AmKRRT5uH30x8dIXDefHxVarM8rnwY5d7ONSwDLRl
UTuABb6AQDhqRLWrcMlkEIOTHRDClWjbOGoJev2V+37YCidT2f94AZ6juS3RIBbx
T6kyeRt64ZXooyxbddjgEvZRvDqWk0xpuN2Sz37Daha137yjPHSmXFJar9k0nS3b
FJg6ob0LYGuVkrelf/4Z7k9U2MrO6PHkQB2o9Vnp3GRarpa7NvzoIDCRy8KeYPnu
dNzxwXoVb0IfXisSDjB/jmgnU6RAfn7hYm5Zt3DBpoIdxv1KiifoMyBOCckTxijq
HrUie2e9/lfaUrcXldiCixeH+2l1/Xq9/QHi7kNym0O8a0gY60OBefsa3Pe0srRn
nNnqeQyrpRKj2xbFoLk6NHwze/kWBV6XfCeVdYsIbxI98GKXr2W8xyMGPpXZC4HE
BW48+LQdboiJJG0XzkoCVZKJPzuxLowTX4qOMJSf6tN0w+9LId05AMBB2AzLhoLl
rfx82ifIVGLeCKuBMiUHk1SbXUZbL4eXDFBZAmjuCT/ldXquk+BfUZJRxIllbb2b
VpF635GMR3kZ7kQC/46YV/2ibwlXYxNYKfAlA6ezmu/xnHocFSntl9pFgWBA8zT1
INeUHOqHfXTdtmJiIz3rEOBVTzoXvuGhyqsFouI4Txv6ZEv13jbDv240z/SNflus
axldhcsAZYWsl0jmdQxi/ZPleHJZocB1FThXUFbJOypUJHxTe2VLB3gfca7DPsCn
L4yATm1JbQDgXNGnrB+pR6QCJgxwwKG1efVVzy8NOIgAYeaLLaPMDWgarMZ0UYTB
6oFo7wcq8iGbgPYGaiiuhyemI6QFuMiUFl/tLl+jC+nes4T/HKFKXWCEzfb7Dc74
gjEbUEtTHuL3jDdFaCd5/EKWmqNH5MABVbbEFitkofSAx20vlmrSvN5KwppGYNBe
gffC9MTtkWxMvShe4LQq1JQjPxmL4G3m9AkEJquZuhEXoF2XlWWs6PhRItqHsyv5
sd/vMO7ojVF55f3CeSKHg7sOtexrBRKE3eW/aSSSbYYxa6XZj9rQjtMFaSLXPWi2
l78g7tmD4Mrps1PT+tONfzf1naXsP2X21qo+NjhF6MICNmj4EvBDqaOyIqz+o3EF
VtfgdWf4glf/XAxacPgRbx8lPwygcL362XYcwzy2C4wy88CuNARFI6K9jouVz98T
duNlnoCojlN3Bn4U5wOrk9dIlulJkhtK+80mb3I9hfCT1AOP4IVdO3Q8YaeYGXFE
R3UERvIj6dgLMaD8S9NOLitmom4jSQxzBdySrzi4F68kKP3k86a/ZtoX7jOjYKN6
0h66/INFrGn8WgoPbZRkWC12D3EMwtC/kGEbt/2culzq0v9BCRjGoTyX8y0p/5Cs
yEnDtKLSjs6lt/A+I4j5EP3knwjHIcgwoM0x+QO7YyqDM3GCSf4RoCk0J3KVXu6T
8/NiOHxOfRILVKCQaEMVY837JCROUKbAehk88pp0Kw79J25x4WQ19Zwf8mR/VYgx
llyyD31s0zmnJCG50P5PNOjcHWKe0ddFwYLRIne4a6TPG5ES+2GdEfdXQbatt+Nr
riWg7O6u1RuPM0+Wy/o3DnQQwX07NKv05NZDddGPAlkr73wn503U1F1i0EBM9t60
SjK9RxbEBqdfy1lPo9IA3QwwdAOndteNHHvEuWiW/xXQ7eCLie2dqYYkVbAJhCB4
ingHu2dGrDJ7DTTEjytqAVkhxCpOEzoGKP4jTlB0BycWFjJrqDJ4c9Ln0eK+zyrQ
vp1xAEzaSHJwl6FnfONS7VaZ5JKdZr0ftqYQAN2C5acvcWNDJG4ytM9TY7hWstt+
lrokWHbkqQ3i/LUUq3N7G6vGqW0YjOBaVmcBwABkioLMR6857xrCrNtlpZtuNW7P
CDIbJlInDveKnPfO7kxYprcknI2mqvcmqQqQ7Iyte0Qvx5uwzTg9WjrwMJFXhfTB
fFxxl53hfIpQSXEQmzQ6b8PiXH7cw9U3YTRmVbbziuBaB/BR1kdwCOeajsyA+MBt
rb25OX3fhciQuCqu2rlhwQY9FleaoYOZx0mHPLn5o4JLIGfCnoqC7kIkEvuskL1V
BHVBLXd9hnuOV27oyeCeXc04dQqN8oNsC0gWcAGKMs+R9ymNiVrzJ3PVPXGVOcIH
XzpLMpVFuvj/ZKquzOmbpeimlnL279P/mHmOcX+RWT9AAJUSLdo56WNz7PvzMEoK
Hc7ivcR4iq+5J6UcuSXa7usRs5CIAYRcI8iKycacaJ5fa/KD2/tEhsSN+vLelohh
VBym0qhNAQt9mdeUO1QOigd/XETbprp5lwqT5uaMFJBRtiFVyVMO0pTvJvUwi1c1
OhpQUnb7J4c3e1sO801TtPJ+RFr8Wl23Nen96TvxXcZRcJBb3hsO+bphLp2AIHjx
HUHeK3TbbSpsFxAOer/VddUUiNrGiE/tJo/EkILFqRNqGY5VGayvZ/yqaZ4UyWRZ
eRCOfNuz/O61A+2dO5OTqlmj4qjR6Rj8fzZqZ6v0PfMk5DVo00gbltDwoTTH34nx
56Do/5iLpaLafRVuAHuk4iSkgSjc1pniDZwuu1+eW49Ut3vCN0urXnOZ/G/NpENX
CrgtiIPQCkwc0Y4D49ebvobkd2LMzC4ho5yyFks0FbQhzNKWwH/TGJQ7FTgMwJc0
QvKWqsMJdAl/dHyK+CL5apw3arcIbIyzDjHL6bVgIydFNdNBqnaHfSSjJeS/6DoQ
9mAivf8AUYgcrwukA9Ur6eR5EGt5omf/1CR+9WEJ6YZZ0WoN72Vzz07Tyk6tFxjy
ib+ExkjBdwkUEjGQWAPVA/ny2ElbipVLiCm1WZil7qz901wGooAVUk4TCl+eI6YE
v40Kxc2/NsubdTcRjTtRynnY+yWHD0czBREcXdqClVZqDWH5JKnim7RcdPA1492o
7AdoYddN1TQ2acI5/McbizGoY/poA4B5ckoguw8NmqMUd1lfGL9dh3x05cE+8I+X
fA/KJ7AxBMpAJhh5VNDkUWEIykaLOfyIVKMe+P17pW6zT+jcopgBm7UZ6vU8TfoC
pJYB6YuvTpqeSoRDsnhUknpLcVVNwgJqSm2Vtzk7SwM9T2YaFlWSr5uk+qKrPg9W
iekNhKhk7xIzESfnhYVly0OPq0fwtbHQfbuzSWNXR15cXnhv1PWvV4H5BxcF7Akg
4WKYyBXLfc9PVe6IuozV0uMHiNVVdPelQBNj6xt3FuIrQiRtJNhe1g2pWsQqICL+
zIdoPUnoJ52Q5S9ex3EWPCQA2XDCEy08Tnkt8QA7qVjaN59DkojPxN4QXUESwvh1
tWGijWoEax4VXiWLIOHX0cEWgIfWPoT5g6jgp0fihA0BT5/kmlYA0fao6+H9096B
Glh4DObmyCShmSAvI8ts+rkw6iUeoeZEGShJNHpMQany10OI4+WSRSt06PxoSpRD
/oscwaB4SFldgODDNHErj5J3jlGAJwmeMZ8/9PNUQzy39/mK5c+pGiHFmfqpYHkm
Dtb+4pm8NYyCy4UqJFAdwq8ENP740HSJ3Unw4xE0hdn9iu9CciKU23gEy/m0qHJp
QIoDvQBqp4ac6//EHZ3adlWXXPUmDSxlkJoCVS4JmyAJRvX8rBZe2hLxJYAcUDpT
21xdRM5CUWoTsi9a50bQ4oCZUgoX2uy90n5lG/8iSf8BdI2KIFWXl7iX4l5FG5wT
0OHm5lJP8uE7mgdXmMGKZ89pPd7VYyMkB7wbfpgeJQ4Mv1MPAS8CUArMj+t9BWF0
uwd/DM1KRaTy0ZdhNZHFFxe2dK7m200e0g/jVzSTssyIVluezoL/3+QMNo2Ui2bW
H4yhVgVZ3PfOSTbKIMOpXF1hNSHpgsKRsL4pFs0AmiMYjGyZs/7lHJXKFpB9ZR+b
tGm5JC9day647QfWq2K2knBSlfJ85rCYtXdj3VSWHh23WWiFHIO9f8Q8nXfn7Sm3
uxNbR+XPbp/rfs+TFJ9+4D3OuTGaVntwh7Yn1AUVpWNo1Oe2iBlI6a0MCm9Yb5ie
CoV9kP57gpcSsTsNhJ3BWcD3Crw0P6+KfBae7eT+R4yeUn0U5JazZCyYOcEzjTi6
ZNrP9gFdEef6/lNP1ikPcVHcXeWtrt7dEiJypKGlzlwk0EYDMiHueYZ1/00m2uMZ
J0O7/3xuxUMJjSH/L4IgKPyMH9un91wYTGrim1mGXUUx6XUNCHDYju//Nrj2jaWg
e1//z0KzYOjrB2CxXIxcqK9hleVupFOoFpKT7Q3tySCWNDLAV70MvZVb0xV42k0k
q6NM+wGHf4RsqSHESYUJv1qFpLDL3fKZH+8Z6RTlMP+XiEIGbxYVhWgSbyzFRswr
IVR5nB65EC9KO1o2uSN/NYQrmZqDsSMhsfe3lFCFBeN3WxOFNiKQdBCovo7HvPAI
eZibb5uix96uBkMl9z9IuYy+79V97CrzImqBjoSZQLLuhSu0pXgyBgzw6JGpYwXZ
pzZTCdbM29J71RVYlSmkqoP+LkvkJXMIV6+09TVZJGFcNkqXqQ4i/n90GckkwP4F
2sh+w1EoL0XNsdbS37qZFqh1Q0k6S8h86WL40BFb62MmTKYm9dfiY8CK90Ncfo+C
QiAb/SMPrgGnVQAmMUof0UPJp4xTPqppKsoiJbDPE9eRaoOI4JTtFrzFbbX6oORc
aNk8YkPoVZKm0T7jDgbj1KDXlGttzo1V7RK7poNOf7uLWZ5be0eQVMUN5uuuYOZ7
TGu65Qv5KAfiAdewE+XNpg6cmncH4zhBU+1RZhT+GsCZIab23aJCOKyGLCmAO0WO
q4tINMmZMVp6b62IQCz9palxIvji+L17AolK3BzJ8wCZWaxr1pkyERGfcjC8/73u
jZhiav8kY95CBk8yFh+Gk3H/HIalHo5phO/IImuWhFeGakl6J5LhO6xtahwLCaYi
6A+Vgf0dNeUQiCeb8aeGd4co9FnjGpe0BwF9+LRkRvtIp+0M72RnAJcqc0t8YVch
oAgxT8Qk8JJ5gl5UiWFPelfnHYamisQQjR/K6/TCMF59sOYlJWnhbvayHUhDwWaS
HAouD5nV59eYoBW8qjPPGwq2TWkBafetvnzga6T/y58WqvCQk/Z7j5kGpukdh0x8
gscrqkzWKO+OirafIRnngJLh2/AaUZ0QLXMiFhP/4R33ByM/ps0KD3N7f6GaiQFY
/U0IoMXW59sdiAMmPAzyVoyeg2aOqlya0mG7AoZIKmApSjUGGUlKs5ZfaA9WuLyD
lyYGHrqw2uQ7OCk8m79NaxhLpiR4aJwafoab1tfidA0AuuxKWb/pMj5Tn7Uz3ZWY
qzpJ41DezkpWnsg73gs43U1Nnbs91TdtCS0TWOBsgvJPhbsxWjSNAzjYEcYn26pz
QsWbMStFy+vlCr8oZvtbiEpFOuhdRKQQbgDC/dSs5nIzdhpa5TeRBZT6WOpxpBHm
hRQY6bkwgkCdikjpTtahrWskx/clnv+04asU/UUrGSmv88SZqmrlNTGwRcP0c1Np
NsVeMhkouv1llb0F6MPGq37+MeWeDqTqwFO6/fKVxjVFgNqn9ZsTaeoXQaS9+xRh
iazSnuTL2ilryTdAbqJjXRgZfBEGNMWxUNdyCHfr4zneJwz9BfmnSGSwjyeQ/b5K
QZSZTS70RFvIhyT5fepJonS1adMHvb49LZR/IAHqV8tpC7/BAwEEpb3hPEdOpgeG
HuU1wk1BerqcV8DOx2821CedXLOSPFtw7Whnw76TX6+OGcxIpqtIhSl85HQBch5F
9+VtUJoeeLQNGLYVkqsy5GMS/wgNoKDUVyOJ4vt/0R51h83v/sSqvz46uLvLTvXQ
cZAA0LzxvjokI1SC5m+Wt8H/n9xuQvwsRiApu1pkD7fX0TFe7d60s1HnoUJ9/zLs
oqBw7tuirnKyzRO8kffOPzVkF3oAmtjX02/6tBrEH7rroPh2dduFP6sjEuADDeyF
Tbws0ag4n+HJ4WDm00rFfnlUMkC9Yhx7sGDIq6UC38stAyy63GuP5KYjNSqeMGnx
FC64MU09QvIs2EbkmkZO60rW67KiST378hpzMTJQGg5F/tvNuF9ar//Dy4tIAoJ5
5QcKMbMVXHN1s6xUC6cq1sexYwCw96hAHprQ+t+Z2GUpVndVcva8qFUbBkkoS2AJ
RtotqIGsMfsLb6n8h20Y1pSKLYe1fe7IVnr8dHvYfC/tCMHvmHaZ3p4o4frC3fNS
Jf3Az4xvHHFJsOhk7YZ/gwEajnEUprct4a1PgryDXdaoDD6dJHVceAEfXAjoijp7
di/dGhpz53jRnvfCqcFrLt7VVgvBeOYLx35xxWGxLXwOI+xkpPPRxhwyfOb/H5NM
8EdTJTg479Fab7nVLVxQwGP7ZAlLCIcaUD6HK7gtebaRY14SEWeBkXNymSORSLrh
Tb3n2/dSBOUHw1bvCpy64nd9t3RYdi2KMunXWCLBD4PAr1JCLhUzc+GiIphyQchk
OpdBbJ1+/nn8jInYuywGQIJyQD/wWaX24mk0J4iMXz7ZXR2bvwOv5wWIzorpWfEx
ZTIcKAtlslvJMQe45Cg650JIBscPldKTnIB9Elx0FQku7zyrwiC614dLp4C8TSmw
QzpKNNZvixaxxIIcFtN9Vys9K03HQABGX5wwrOgMmWLPTsR6FRP7AzFwTKYpvmbe
NLKjvgoOm8FEDVK+Im3PtG3XHADZ2MFul6sma2XGM70XG1VRbIv0UyvSIEUxywmm
4xAI4U6h9JFibC3Ki9spJQwRmG/7SSjxNY8BAfA+NYj72W+MJySUiaYPVIRo294n
19GYwaWhBeaRqZfWRGpQQSQjd5kEgC6B0ynO8jRf2bpTusyhkUG6qUveudOGkvr/
prEMRBJYiFFGfCNlJ3XjLVRMrbDRxhnRYpn0sWhXzh3f1acLl59X8OS3ydTpXxTg
7y+nsjqpPV5xXuf2bOZste3JaEfC/ZrqPp3emA+4+505lxIrrlxvOUBN3Rl7+//8
mZVb8cfPO6oRwiNtHwm2VsAXOHClEvDazPQrex1181Ory4GZLvNiuNidQm2qg0su
0RDjNrk/v+W6SVrX/Z6hb5OQxqGzOGL5JisD3fnUcFLxOdlgrOSfj7IHlOpCQUlv
ku9QdvxrFEw7uF1hKkKBmVpzWOdykWsdnGcdmF63IVakIrQ9UPWkQtyJSzVtsLgf
xzaRpWKaSo23xr4gf1GzVYbY/xg7giXPS/ltggh/DIwEgIKe1Re1jmmP0TPfm7Px
9XigZ6BKquSBRCqG0npnnpI/wVnU7oPXN90WXb77yTMubzc4kbUjCvcwk0Gstzhr
LO2t6E7XUac7Nw7s1W8ey/xc7iF6qpIz7ePJ4rAYh+K4X7mfGObNDqS9EohsYpDt
w0hSNZX0pqAGN2pa0ewZNwUyYGIWdxVxCo4Qj2qz5ZvF5iDtyT+ZBMQ4fQt90seq
vXlKYta4eQHkzKnG4LxOJB0d3a4Ah7aTGODD5PDZqiF9T1aZhScRLIWzf/oMyVL6
murakUW5g9pt09RW8VexvfcMWlvkymXWQi4a/xA09Pmdwzt4u6v6qFpRp/ffouAm
9l6nzgUmbyEo5Dt2EdChC4M8lc2ElGY/865Syc32aFVRq2dch1fjsGZCZYqKQqjb
sXydXq3Dg3kezTSLSrwuUaBwVL4MJ+Xx+FPTaawNYPiscar0tpJddEoWd7Bwbcex
Qg+Lk0T9drKOnUWlOiABpkkh2X6b/RC6miz6TNkuxZtAApfJ8N15D6Iwjaft9ykD
SPjUpC9DqcQZied7VK3N5Z0IbWkoFk5GjsfrB36BQX+Bwrl4CUejVDKsdnoatLta
OjOtEbQZlhkbw7XubOOrmrE0lIgPePSP31m5yzEWEeT8rnGZ/v98KGobcAyzQoyn
ELp2Hh23QHMV5GK+IoUeehmUPbaX5RqDrWZWqj5qv8c2RUaDEkCY0AV1DP1OnXSl
I9ig1kgmU18JRsPv9ERYohaD8xCykoweD+xzVP3C6/GN/fJE463qoOgOkqYH69N0
2xVxPWeMMjZt9Fz/MavZ23EiZYFo76TKrzPOCC3ZBrG2JhzMs18O/4gcmT0RxDsr
QkxaNRtRe3FB8r+VxL3tkjpHsxBfLr7xu2f6OZwuIXxQEr4UiznDYDcUhs5PaGiT
VwPlofev6szbbE4rKFZPxiKfYpm9nBTNrQJs/rq2Vbk4NVcwupRLuBqSjEVwYKsd
40uNYVZ0tSapD71gj+2sebxUe32A+uJ5WVPLr+yQUa3ljv4D1FOFGCQI7nj3i6HX
Hx3KQ9W6N0TWZo0wFJMHEwn4cfwVJ4g+FRJVHqSnaoYjc0GVQUAkTvglw63MqOMj
5O/Mkr+BdJTs4Z+hR1bO6HrYKyX8Jsu+yEKySvYY8YGS8+gqwBZwo5Yx59W5LZt5
C1JsZ5WuWtebXxn2d53M6AFhzir6Nqtt5FGuU7jgJA9LzkFzBfHFEZrWHLu1mmzL
OduiIN3Rjar1CC0d4yO7vw9smcxs5PRlcAy3SJ5srCV71Un2uynWHMXNm1GwAbIo
LP4LvY7X7MIQlmuteuPxHZ77dKWx+2eAzNmgU+iR2AQi7hHLQOCAIJTuik8PVpDc
xX6Qt6tiI/Su+pXHAI1iALJmdJkA1GrX/cXktjS+MZRrl+njqd4bTrgc84xQS2iq
iEDHOVoK2favUHf2PWAUYHPFi1zIBfPf6PBx7ecWZmwd8SWZUEP0QJnObN6HR6pZ
G9psvuc+rh/13Wf4eyettztRGArNxaEFZgB87aZnN1flOi1wv16Z70rKPSbsgjan
M/Yt2EQluB/3op7JLoP0DQWjBX209X+QtmNoO+ezFdk9Ndqd/znNB7XWtoMvxyAu
R04TeYf2/Na1VThTjpqNCKnvhyV0i0GzI8mugsdAhAFM8zInngCJMuQGPBg8cSq2
6Ssi1kXscmdAcAmSRPksjcvJrC2qyPudi6q1QcUR8Pjcc/gyhvMCApsqGdUVWoZx
nawSdgDIituU9piTbJrPmPwfOkKH0k9S3BYY5k1pSqVS34K+zYgD0vrgFQH/KPRG
JaG/ExrWviEtgGXutSLl80NBm2slhBtZap4BYkRQ/ewipwNr7rjR0U0CBX1aHAio
mHW1CyKH9gctNPqLMMGKp86vci3DWgsWVJKGVycSY58oKzpJXjaz8i2c+OvKRF4e
m8ZthUQhDM3AFuroqvuan/MD/t9dI51/n0p96vVYdShGnAfhBxQoyhGP365d7jWl
MENZYmOF3owsD9HW1UPK+gqGf54UITciO+2aveakX7P98I+8OA4Aa7wmpGqrKRLQ
bC7uC/X4xNJMMaipdndwlfgc7/qWCB6l4Ef8savaAaK83sEuzOMA/jFXyqQ97F15
ZJXWc2DiaKMGUFzT5+4nbLYrKZtuuQF/Y087LMVLHWrSmkrc68sVLzPj05TnhR80
ZjPGRMFil274jQ9E1ud//tFFrjBirh5z+nEJ0wsdR+7QZFvG++n8QFcXd9VsV4Oe
achqegCcaP+AbnYR/Q4zc5VDXjUQUuHQVH64XhmYQt7n2I+1Pws9Gsnn5ZMOglEG
sdsnkwwHnU4jtyqK6eB1P2nYcuZcC8L3jhbgdYBB4sQO9ftT46Mo1b27KWjPOkXn
JeYnp3t0nUVXD5p2Lr1ZR1EordmPegEeN3nKQoM/gN4qx1GFSgz0yUcc9M9yXXGQ
jPWCRQM+lXpFL09sN5dK74b/NWUt9vFsvyGABXQ5vKbP9KxRCTMyNDzEACTVBmOd
ExC8Emva2WLLfn5j526w9ypfrihTXAEYirsM8RqI1Y6jWLxI7XMYBa8O2QHyPNfh
4LB88VckcTdtamU104cK014KHRlSuG180vf04tbSl6YG4RMz/U4gd/84HUsWm3X2
93eZH7H8uxxCKe0z7+Manff9zRCf8jD4JK37ppyCaAPfSlD3WNGSQcP8tqqXuRrb
a9YJgY7NRo1GkPkpLCkRdQNeTQ1NCvPspnOYRONLTFRDTiIfds064OfaIfPK3OXA
nfWKyIUk314c8NKuTeea1kOg10kp4P7tCHZLLNHMl7elwa0rYStKASHMDO/SHWzM
MHWiSBrHaEAvs9U1SClTZNCrsf4J0yvfzbnjXU7yLUMsKdBXnNHrQbEyiz44hd9A
KzdpWs0ro5Tc6m6H+P3dWQkH5Kxa9Uk+WJ5gGNxDwNqT+zPeuaEdEjR0so03Ki4o
pxub0+b6Z1RPb0zJSrylvtk3tR079binwk3th7INiWY/bsS5NDDV8SyJX7WFvFTO
UMWb9vmH2nS64FvxNXAuVU5KGuJx8GE/4PoexiKYsmDQ8uhW7mgA2XnKOC4WKmbe
1dJrXZFGQ5jrlceR5WqdZFy6TTSTGiCcHR432t6ErJbYfteKsNgZC91fKXY9BZgI
bgHDLIw8cozr+9uFTW3XntrlgqPZM61YWifaESQ4E3FDwnEBvJzmvMtN8niX6EMm
qVdlHITelNAGcTY8uDkFbT7NTQgVej7Uz1yXEuOCKkmpscc8EXztx97dQCL5c/u4
i8sTspkkUpr3MXwcQzQKYfGA8TIITFDDQJWSiXmE93Omjp8ItdldMk4vBE6lVdH5
wMVhXv7V/WqDXO67jXQm+LfDXzPCK+SzJerJ3L9TBnSz+Bo/VPUKYLPY5bqMygT8
h3zXVkgtFYrUK/H1T0ZNO4ewlLvwhlVNzxrTJxkmrPHIBKm4ji7f0bwGXum6fjmb
i9rd8QJ5FpNqlzzPdgdR4h/Z26BL+9qqYIlGtXBKiR6hFVghUeP9UXy2uxWBYjd6
+O7p4aU7bDfZ8QHw2PZfQ7u369LCZbqdp7mwZM16L4s6AiHYdN7Z5yQ/Zi3xqloF
SDBFe0exnGKjI+QGaKXo2TKIgvSm4Qm1puNZ+CIqSYMvtZ8mOCjV9ugi4/O7pfH4
zMinIALiYDs0TUvisLdz822RJf0DI62a4gn132/Fs6RA3AF71qb5jOXGKFQV+GXR
0EAiCs+swq2+q2WRU0GnUpvyI40amDNKqvlIGYFAs+0+AI3a4hD4ZhTXB5Qdbxwc
fHl0ShtoQzK2DpIcY/7Nl+AjIlHsG/hpUO16LjikhptQCwkxLv5jyh4Q0NBtp+Q5
CzOTnzQKSFJ/lAisjdX6q9+uCdSNEyvTy4HDMg2yenBJTnNoJ6HfN18oDwurtkSS
iFJmFtg7UHsIw1LTAhLw+BlHP87kDHTjwKIMFVJ4tKPu75Yvsn44WcXSfSluuehP
mQEAzgYXUll/lNeEsUKCaBIIoYxP5JDh5NzgqA/Ve9gidKpEq6VC4tAtcYSwQ1at
J3lBNBaF7PDzI1LCQJOxd/IafVdJ+mL3xK7mbxHNfBU4BflANM2xgmu5lGZIwuU+
xhcakEozuMAFPQNTP8esgfvRepBZUJHTECgY9HPIsi88kOOyRIwIOj4gIoFD7sjw
r0ozHjpQBwxwQBR/9kkZ6b+UlzdatJmtbziJHmg5z18RNrkglNLMSYMlWZ5lH0BD
Bpmdi+dv+xf/s0WGzl7t+38MpmNjg+Estlbw5lMZ9bZkOk7EhpUJOGgr8Y4cjDQ1
dCqVV/ZGftce+TNygTuACrQtImPbCcr1hTH5RuxCvvv+CVrCWugYyVi65jQIYnlo
v7VSFXBg3lIjsqjMDQRt7W/g32JgBccUSH9drEsi2lsUZiFKNzSWX6YE8meQf6cF
UpcRZsWUiqJaJQ/z9OpZqXZI9OMaJ6LEHV7m5W/l47Kd5cEKopP7Xg12L3I1sg1y
R8V+1cxyTTPwO6TDoXingXKACaJ715JHgk3V0Gx8FLBzIzR1MOKBnqD8x8TVEd6Y
8sJT678qwWr0rAOCPXZWw+bMAqEgoi6rSM+OutCqpDjmpOvRcdnLz2gqB1qR+sqo
MM4r4vTiieuNS3mifRrPBBazMy5EW3ZSdT0B4fB06F1r5Hu+QqmqKm/4wlFhF/7O
WWAXdhWDSAykjKhpT3zPiyQXpO5JRiSWYx9gJzdL8azl44ce3Ip123ru/BKpF8ZH
UwdKgTIEzfBFIDIAteGIBJyF37Finbvbhp/PMh2/BMYn0PY03fOwQdivYsBEbqVo
mQ+dbn9hcYg/HIudHKm5AwCenaoTAiH7pQCL5CYfLliqbKxy5aH76LKlhAqyeBWo
illIcgNCAbwHBoSS1KMsIoT4femtVzilutT9o5S05Mk86K+iGdz0jAnZkF5Zm6rt
GCtKoLz/cT/czUAuIS0TE79Z54NmpuCm/xjDIl2RPQ53zBFK6JpcbO1t70keFRAV
hZ7nTAlAe4nd4zpcyTCVXH96jP38e6xHwlFXt57n897hwj5bzYgNlvtvinO5TXWH
UrbwLZEDrDdneH2ug76mZcsgpvQWO+J0PczBjlnVsRNa31dxg6dkUCADXyj3gvhA
ZMCkSwJUnFC1HqTiBMWD7ZFFZPC6uFgVWOSorhhC05chXETCbeGNdDTB9Mob+D1L
l5FPyQBlcU/sR6r0AWdlCxbKZ0xx/F3Fplbmxk6BxbqnnQxp9XDa0i4hWooSigLO
OA21Fn0j7HXjeHhU/oudYrNKpTLV6y9p3bO+i1cMEERnTuo4rKWdrGwH16dxQ5mi
/0x8QM8EWIG76YFv/WGbDE2Gg51KHVQ+6RV3kO28+9dwLHrSHkyy/c2pgtN3nxJ4
UNpSvhdXBLURiyw/IMfI9n8oa53DLiRWyu0PXsxgrFwu+sjPRWS6KMi2HZqPtoNb
KFtwU8O+pcGMz8LgmyxawAzgqs9bJQQKB5ut/IO4N3rhCeNUhBsMHl99yKtRf6pv
z22N+Y9FRnPMCeKU4Ce/3p5pqSvUcHg5BOFmg9OzRupCuLClZ0tPofnOufpSleXy
S2IG4sL3TkRgH7OeGLYtSNIggALAfacmL8vCBIqh741uhA1NYczzJIvsKIc6RoQt
wQQ9Xd9OWMdT3WcmIfVaOzWA6DH+EnjvI7klfkwOlN0mx04N1ZhNOHVaskYwjKiT
8rdz9Kyy78Llqe3dMmT3pSK9MsU7C2QYGUCYddOQj8WAXRX/nW8GHrfTaPsAMbe4
DpIFEdhr+oneChYjCAtd01OLFAbLVutJZMo/o9g6JXAnqRInNNjbRp35hfIYZx4S
iSq72/CIwTKvbPfmmA1FKtXe4CqSjkdxgE95IsFrocF88Xe3dwiYmDd6mzo1TBEg
+xlA0Et9t6bL8VAPGw3Hswy1TmV+1am65dpzprkusa3mfrRQMUQBksSi1T9aad5J
/6zYn3ZuQ6/v9i+budxyapbJAPofPfx+L3b3oeiAuzLjDx2sYO1ikzu+fF/mmJwg
aOy/9DTcfhcgjzT+D7NOimVJxKlxJ0SgkauSunos1OTop07PRFHQabbIoE1ExWxn
Fs3BSgRuiRuZWt2t8VnALffHDI2pLtM8GJPkYDSUBWIdXTwjKdOnF09eymSxcXRX
vtoUGHyZ09aCDmij74dCjlp5SYbtV5lD8NWMZLBApbiQiQDMY8C9efhFG2Erz588
l+MVKW1MXh9onkdCOHXzOr+boNb1yQm/n8uGvhWmr7Yw9Lr6x6jGMRFkpD7CYv2p
CPNNVws7Bf+9EylYXHjLhIdIvUpdiWl5urgS/dA7V9yR2pny0bWpRr61zdNcu0wa
ZPz1hbugRawo7wMbRUniE7Z9CUd8yifI/69lpTy1yye62AfJRBgEhUAnuEL+wKDm
1jKw0sxD56Gq4rxxYq3ffZFMgDOGuGhD+drZtA2ArTuLrcycaMTXmfGKZMAaNVwd
w3HXwKa9S8BFxzbEB5beyPv2geIxczn2wV5a0LJPzAkMucbfLNSATokf1Gb+vnTx
sqiLYfNVbK91OsIl0fwX+Wd99NHuSmMWW35UBv6c4l3k2MleXxIg/eYWg2T8LtU4
ZccSqaMniY3EgjdhJswLE3TG6DUogeY3d+52qICcF5P/4NYU4f9LWnRl1qeW0o2A
OqHB+gKoKpxPAaj8xFzQQ6B4kJ5IlFf+Cwn7NmiZCPQenw6wcRFui6nteTFW1J3i
wG6lVwdMc1BxgCDxK8t6W5896OCk3WVF2eHB7SLeHYIcfYM9SO/8iP7l7ksuverC
pRsjLEvZFxK00tATuaC6l9ws4zVchd6px8aIqcyt0vno0VVDM5RgK7ADfhjBfsTH
DSX6vB4TYC0ssnX3x0tW48iIjW6IjLhI8YMm1VvwSUzMwkceAx7e/Ml0X4KNpRwE
BnOqCH12y/f/VEOz+xVgL14zQD4mupbyh+DMuciBhRJ/YbSAmWazulyIRNVTbFWC
qTylN73AtH2pXaVXUtLYNFhIkvrJHFucqpfB2dfkb4eR0X1G/GzpWQzIbVHsE9Fv
wwxWRAWBu01sgoZDOvjGVrcB4Bj3NFAK7NTnj4jy2omLnQHkxUVLx6HntM6gpzw+
ut8UVvzou7IMb+7m1to7Iib4dwJwWgwh4VGHdG0CHDoCT9G7BIx4lhcYnFvApbRr
/krP6wTCfCsv+txDb2VgLjoXHMLyQiTf13aEVV2BNijnJ+gEBRLnU74eD/vq8RDg
yIpleW5bf79t2dhkZhH+a4sks17EDMKjuSu/OpE90pmzxuhmguqaAb7fFnYlpvgc
63QkTdzlY7Nmv4+oPlg5g+Fdrg+zQPKXrHtCEPykSQjF5Ys+3UyCJvi0XRwJgrOf
tfF+KIFblqN0N5+TgktZg0yDxf9R9YJAHXh6tO76g5Gj9fgmN983R6cC+JVs2Awa
TgqiCaV/VCTSBxQSwFw5DnKd1n5ZBQZLILkDVakbPv1V+tj+hzItMMnVUu40VtIN
kZrGjzqefRu8ZxXbGZovVE+4iuYyDjqDqRAio40zUM4iIvzrgQ4ZHshij1LnzAQ0
iZTp5rn1oIX+9DlSfYZJnfe9Tqs4MMzfNfBaYr7QxxWo9r+uYMga1I+2hVE+BwOg
4jC9rfAJ57Th+o69sql2o64Jyc/Q52fe323PA/0KGJ8C4wDTcWh8p2SYUu4FMBQB
PC+BwsVl8NxtjEFo/Xlv7EdwUXyxsYIU/Psn557CgAweDYc01JN1neCxqD4wcx6b
ERT4nV8zP46s1FXP6hrJ/d8vlu84XP86y6c4kRi/KY9qgkRaw1fV6y13GMjpvbFC
jQqIpoYIJAQCTofsyHCU6MWU1PxhPed+OpAppQb+vE2gyIeaAD/mrL6764sjfUdI
6wHG0UH5ZYmfsbJlQUb9hUNzgeu6IZoIXsAvpIcgCdTnRmmnJGFpBCFacOufWeWU
QZNo11SuY2Ws8/kZ6sZREM3eof6H/2gjcLUA1pGCqJ4u6KAhdqxGfVAKeU3qCmZk
z0u5aL1cV2BS+k4s5oQqL9EN/9iEGhNsb4yocMDiPAWwbkPHML+/seMUDec22ZtF
oq1ZOPbjgYsKGSnb4p3a5UQefs+vwGlIOST/AuNqwIa66tSu8Q1u6Drco4sliteN
020mNoPd2yNALXo6Pj05l21Uf7xdVifPHAS0s9ftavjrxIBDcDEeDnJkaK/EQA25
IuA42FWKai6pj6msx897pxzM75XuYijwBKyuWj239Y+oyPz/HT1t0BUTh/MXGogH
UaEhr6Hcp3ISJsqBD5yGcWgpBNV8PkFOD4ytSiOghmlKJb91XugX5KcWMj33yjAR
k3cTeweLkmwodSzW/2g5DYVu0wzRDwEOvHHJa/hmC8lAHntsFjLxktJ/l250PUiJ
im/DUKZjCirvSvBGczdhyyxHODSHymKp9x6SV+nJ0cnpEDCgpQ4PZWpg4gDuHGlW
9xvNS6tunX1qfwTAOCywfzXHT+Pl+7Ihg/7yKKbYeEEJ6Cwh0GUBE7NdLCg6TPX/
Tf6rBLVTewcQa3GmeotNl2LxusNjKeiGRPGb7KtTUYYsZh4JVXBO+Rz5R2NEE6xW
yF4UyAV04hrMqSWl/9LnLYZKfMRvaOn9SUrmBLgp4VZ0cxm6fzI0W9ei7EiHqeNr
5vfw2c5k17KkAgXTlRGZ5Wt/Kf+jKORJJ6FKTmdZgeiq04EMirDidl/+huGooObs
6psUU2LxFxYiBRy5I7t1U/Nile3wVWLxDW9WMQqF/1AkdRRWa1iQzIREDiwqp/km
6zdUJDx5FtlocLYQLMEujc/QuJSZNwGwDdadeMOmyqvwp8Vbt49n+eHaNco8qePW
F28ijGUTaPmissXgDVqDY1iWf+j7j25zulD9a7v/WIz0eODlyyykGlfCgcLY0oLH
D/QDXjv+zq3cKH2SszfKC+2B03jJbCDSwAxPwv0fB4Zj9k9SA8mQH0ob1PNZKEwt
XHM4zSDIb+hpgNiIuaEx98ZWPS/bXIJSHsTPNddkiTu37j6NgMuQeV2MNY9l4xMq
GM9sa764MzC1ijqoXpMFACrHtg/cG8P3h+bD53u00F51uby7FPvlsPdW8KTBWsBH
AYHJq3FmilqZb7bCqUlhpViB/X8eM06vqUVq+agjs9ThayyZRQ9TIJP3pKmCjnzN
lFC/GktjNjixF2mP5nuotI7kGUTP06O+RSdmKzYjomMIBLFGg9tgeDsovFs1lOu1
+LKQ7QlyqkM2a1cjfenVBHW6H2X23CJgOws1WsrQW3xOBQje4DjRYolroRpC47Yj
ENbS9J+mYXbv28ml/wOAQdqXdrgAy57Ym4mbx7Ttw3vFpjQaXapdK6bOlAX+TOJE
fB9vgdLRG3hKkt+0HJCq3HvuWE7uKLc2FPezn5/FIeIwRgAfTRGJN+QLYHZGTeh6
7D4O921g6BiwzoeW3Ae0n2hkfP7yC4AuvHHBWLUbwsNq1iD3T1Q3cDlzdgnFJv5D
GEjzlFikJCPrG8lx5ahUrwxhxgQGdDb9VFJQSGpuGbv3POVtUsLzhmkPAqVJhz1G
K1LkLvdoyrSOtQtR6NWPMvf2v78lrA8tRA2M+hX4gYGw5UykxGukbJNM3O9h/S0u
G+TI7lDrsyjf7RZU2QVrRaIbmfde1I8YLC5nILq3+ihvVNMmVIheonn8pZoEfdlp
fQGNIlFZOLR+2dddqJ6+3TYNxrQFy3ZdAi2b8cILvlGb2GUfm5UOAMEpXFSKT+qz
JMhDUJVgSe5W8Ip9hTjS7dGArQhObGbKBHP0zJu0rO5+dUnSUU/uijFWPtYwoMl6
qCC/zn6Nd3ALyM7NSoVWdXBIzvifT7dkeZ5Pj2lo6HxXRmsgWcZGhlJN86iu3gq7
EGjYrl+7HVq8wka+V7R3aCkCLGmFGFeYpweub87NJ9HLaJVN0QtzTWSroWLBz/8c
K4T/gRPEpkiuUYHziabB/bMKw9SNUxY6WA/Ayb3NqXmft2eEVVfh2ol2h0KPINZH
R52+U3PmOK0kWxBBgrDADt7QCDeW+GbgFsCccmM4KAoYnpOampLAQoDj2bOCTPv6
M9ZlZ0kChxlhn/sOJNbA/W3zS51nf/XRIIcRiGzrvAR/eLLigfaS60lJXenWFP3J
mV2cRxct8Sd8Rf/LbRhwnf68VKrLugWRYocC5WyLH0BJnlf9u5DlAeJCX+0k7JcW
lTMiAHQOwDXaoyJZjnryWr4c6ZgDcYS2zG/tJHSUETAusHNUFe6evWB/tqJkjl78
T4xSEOn1ld78lbZb0FN1pvyMZeU9a26Dv52b55aqiaQCW8uL7w+7Er4EILqrP7y5
byYKMabIuRWUu4JUygp2/wPOQBxLP/hiSFW6cIoj9ZUVsduBUsbXkmuoEI5guqnZ
w/gpSOe6sWJvJnztDyxc+zKcrurM2SUh8y8P7suW9Nu76ZK8kYfjNnlcFJT2QvIV
+dX5qfjiYEsCPmHc8L4+WDLyMwR2Utfrxp+h54OfssVrvAf1L/JmMYH3SM84P5iq
51RiYZqD/LCD3wqgQvRpWn1h/2V5Czd3D/DQigtw0R6s+ICzEVcujSjAR4B6Hz5R
iYyoxj0D4rveYaNmye3AzzUxluvgH3cHP1k8yTEBzQYHxTCfHZQIHCZl57inBFjB
WsxXdEvd3OnwhJc+xOHT/sVBOjBPlsPZS7C8rGK5j9Z9KSh3jtO5rbFon0VRDlqQ
y0FyBthGrzyro+/HZX9c42skXmiZqr75zAbtTcKr6D4+fRuPPALvvcbCqecuWj58
9dAr/+uTt/u6/1x30UsqOjcmsw8Hk8+Lweo7MXpEaJmOqMssQ3ePVSQJM3P9fG+M
ErJIxan/QfYlUJvmKs6tWbgCnFvgCJyX8EgHJ2TutTgj09zh9YONobKG92qSe6gZ
BCWnakVNUKZi/u06yi54zkXWs+vVeEedQq7Ib2ntzZZYBpxw+G9uDCTN4AkpcLu8
bGap89aYlARuaBT6hj6Jtly4mIP9LlCyLxzmnQfEMFw2oyDIkz4pGKfhUssxgVuc
vIFiAspi93jZ2rN3uUACKgq9jhQo309cjF0An8wN6CBLumfYjD1/l6OWTs8G+U+F
drek3A8szrlKrFkAXDvFbN+fjNzVsnhdKdeLG4UyzwrL1pPRukNFx7a6V/7Mrac+
5pcGmD2tzPcLqeooDTANDqnLOERYbG5smiFBXzSm3A6ybtljpFZ/dzW0b+K0URZA
iJUvtugEnPkwymP0wyhcKSz5CMl1WNDyuThNpOzAgxTinN7LJA658he455mYpIRa
C80Wbmt/NDJ/cAphU22YPsVYctQ7jHZaxYVba+mY85gxqA43hMm/iTUUVLVPt5T2
6vCDzKrISzof5/cwYQDtJuEZ1cyAmlmB9h4OFoF4eVSyUMvvCD8ctz5bbX8MGDHh
8x3Gu4KwY/pTWJ5752/DFRNaDbBeNoaUwQDyir0z7tvLM9bCEqZKH4wpP6p7gLAw
Q530lgtbbiniV6LcegyQUaGxKRlcDXI6IZReRLjvi90M7AuIXZcVJ+8vTkLQiHke
hNbjY3tSZv+pg+bU6+xRJbygJA16Y8IB/TNmm5+N9O3CP1YeSYlwYqavgDZmdyX5
RphQ92Pyt2CxaJTwadyVvUd81iB3VjHwn72QKcTTuKylifTi/dknP/qP9xQ9owVh
rM0ZFgSaGWr8S4TJv+88ZvgkyZBcok0cg9XKajN0DJmSwJKdJeCaP7SUc9XoBP2W
DLiSZ1jRH+wHFmD+ZSKkZgo9YLvAjZ1PmITVgMdIMlg8+bu4NIgOLwLqaSZAGEvw
pES/HYi8ZLguiAnUswa7Ntwth8XzkygSJfOa1eCciS8HkooblXW5FX/W/R6iEs+j
QhgmVMDHmTsP4B8tBExxcRqpRUOpGjp62Yr5fJ769yG/YK6suJTDlSMLVjsLeSUn
Y+ipAKxCAF8afbShtUQriDDDivQ3HUgcTGZ4nkjtFRQcqswDSP4m9giq12Ga1DPq
WN3/daBEPoJwrCqUX0u6kPiS/JwwC0hNYTu42yTzIrpHAnvwJ4xiscP6hYrcF4ZZ
ku2jejpvcyj/2fYsKKC63Ws20h0xhAzjqaaOaRKR93P5oWmRRoEUpLlsUTycB1Zf
wdP5isRXXzfcRdLAwonoArBRI7KN1ElFDeT2PD19tgK7eY66YHXEFLvHWojTBk2N
rJUtHXN0P2KJkMxUCdZdMmFPY5zz0x6PpSgC9wXXLALqIQpcl0b2a9kQuNRUCUVL
+h9YACZmj7NWQue5j8vKYbiwBcd8+ywfxG6HNhi+BORXFaff0V9vioCC+/+N6oUG
QfOrU5oH9Xh6/foEK7AbvyQhroTFYV7kmhDiutmi99B0mOVcm8ZabD9Kq+IMMeiy
4dRUC42uVsa9i2+y6LoWidUkdO3WHNVssvY4uRdMSDiLg0XjzTXyLVRfwwmvFlGb
FjclYBUwVuz/EOB1eEsXgwKq36aCgk15Td4F/mn/vs5bhLwq9NlFnhhI+iqHwnlb
HpsJZMEda4i611Iv0xyWZDYOxYNWNrqnlO2HJ+B44IG+bAfBAEsi4tJpZ/wufthU
F4k5U+tdd3bh6osYSWWvY2rW9su3SOn1vWZ/2GLHwarGlmyMkPcI0u7sS1uE6RS3
LH5frlhLr2fTnoaRXSXQZ0/uYRpP1whru1rEIGuEg6ptWWgYybv+tG9KK5vTG/fn
C/NFC3i8lPM5HUuZOML/iuqrEvn3P7hwrz/T69pgZlHXMzspPr2oZy9O8VDhgmnK
cJelvAU7boUDd8heQrxxgFy6T2OsWBWKvfpmMi2ypbKzKsyxwbxrzyiluJwfpA4w
UqMxgxsa8leGbZMogKLF/elnLSlF2ujV4B+r3yCAvU9gjRxBVp0xrvjsLy6DVq8H
YEvrMr19+Fx8x8BY4TEZu6/yL7DthaXnFh4L5cOzmwS7DxSmpOUwqtO/ycXbw5lP
YiekscwMqJRQLQab2d8d2HO8AO/SX77AhYfxFYuHjBX8mAhHWgoybbfLQAtw8PYT
E/NUKAIJYDC1gUiXFc/sbYPvdAxE+ZTJemGTOQIhIeDh1PHugkNVC8rbsY0ompXM
OLwYq+pGVn6lLO4LNC4qDiZY6mswTphBquntn+udoK3Bxb3SxGQeg0xXlAsWvnqz
KBjS7QmcfRergbwaMIa96GomPQ4AmfkYb6oqffWVClr27itgqcidGoCKlHdewE87
4IhwFWbEF/GCXslvINaFmqPh/qnENUFkHv1ErxvU+q5XZ0Zyl+p61wYd/tkrkPkV
w0gFkiMDPSkZkYt1JCqIHz/UdIbBXhKgfb7fFmySHDeBIywbBvBMiuc5ngLic2PH
GwnILBi0pUlg+MWOJg/yk/cB/jcNfECcuXXifmmObulyCK9Xdd5n342TO6pdBvQr
5JRUerbvW5s3Zlw00jXqkkVjDWdJhurYJUK75h1s9KlFCZT52IME3lYrMaXq+B5Y
2onSuCYJiYjh2M8ywWNTN2bsLKAG3RzMl2oNRdmOQiGquE6YBCohvx44A2D5SPNT
xezFebEVjuyoYyaisFeAaI5WgVIqWMPFFvXCMxyWcOnnESTBVy91lGtBJ61RzJKe
3V0cD1lPY5EmdY53Vh5tZjRELxBuhe6698v4/nFDsZwOmkyJuP+1U2d1hMqOJixB
DYU2zlNtE0GS4Ww81+GFEMgeaGR+NU7qP8vcx2XfSRbDndfDuiMXl5TWm1WxbFlT
rIqk0Xr6iSRHQrWZWj6KdoOzskgDf0Mg3nZOBM/ruHq5VAG60m4Sga3KgruhkeZq
EzfamonS/bZ2wIpHZHhjEEVbCBQLwYA56gLe9rLI95M6fbl6M873XGPKd8HrEHKo
MNGmx8NsWhwEV0z37korjTp+z5HhoiTgzy70enwKO6RidRX47xyhaIpKuPQDRZuL
vmsNCJW0pnQyyorW2RX9n3on06Vh1H22LqznbITBFheq8KU/kusXMrAfK2AIaR0q
MOv6ra7uB0UTPOibtylZ4W6515w5EV22jY1+nrpsF4h1HfaiEldo/FjVGBADB+FG
+ZwtMIqJ9cr5fAyoA2eRs3aS7pVRsZ1t4rKaEyQakK4lpq2w83k41XcteiFSIqWF
exqOMKxEfpo3I8QB6MtxyKZmUAEkvQFSWVLUnmLw2MA7FfCZGhZS2weGAUBQj57y
ECbxvXDIcCL+2YrM6/oFEOZ5yAHU0NVfLEaPqYWp+w/u8gPaZ/pzBNWYVZMZW7Wf
Gzmh1srjlILDNRnNtEiAV4fc1A9l2UkCRqtyqBHG3uHdGeJq+xVuSSneWggcasU1
/N6QrYzwpeInW1dX2eCQ1uo0CqY67z0eRghi/vxzZC45f9Vugivbsc9kWcNnuRUK
VdBY39d9sGYXSTW/JZvJ1nXvzsTjYM4t6QAPaNuKI5u+KLsXrwSxW5yiuX4+VTC0
tVkq/UxEe/JS1e5oAO5rRlWUCfDNjquTkqrzNCClF36vnqMy0VcV1QCQLBbi7H71
wGiZ6fmmESXi9K7zDiDhSIt2q/QEOXJcIHUxyEOT2yKDlmrhRcA8XlwEDGmf7Y1U
/49wzb6ERHT+uN13o6Uvj/V6+vpgbvNMKe0tJG7eyKL/sVoMJgygnmHE2YR5kTo0
Y2l5UtHgbarQ09QcnOu4Dr+Dqbysoq3q2kqhk61ag2hoK/fRZ9pUf27lcOux12aD
1tvxyeKmnRBBDPqXQIDFUS9aykKC0Ddi+UoZuWctEmQpJTNvbhiQ+Eo8GignGT/l
DX0kaAareKh+S1XObHpVyMTEoY2jNQJDASGBY1a5vL0q6c7cfaQE6OTdXbDvPsd7
NMT2Fhe4l4Lh9SIXpcBGGHURSWGipxm+cw1RrA2+2UAw2aBKhdJ2l/pKNhFo5QUt
RVFhep+gC4H5TPSUNcP/ElBcjUljXzv+QGZJ87nonPxaIioyefYyAiuommtJNbzC
epv/v8YzU+KJZhxU0F5g7hbxusK1jYHNcJ2J74UQ5qcqRFhOC1R0aI/RWiToFoQY
VoXC9ayOc/Deemb/Sz+oI6yGZSINOzoeEcPHWnu8msIzGO1BwwIVSd8ElEQN7Eit
n8BORN94rA5ZqNvLzQwQRdkr4VhN/zn5EXJINQKDxKBkJs1fXFtyDm6Ed2eK6kz7
+UAgsTjAxS2jgMB/meD4605QWmHtUZnD4e56dC6MNWeNoOQAJtZF+7gH8SoP2mdi
+tBSaMDBr2t+/AH9i4gd3YTg1ivO+QvML7vY6dEO8Y2zMcFI2u5n6LgET8buLy7l
mBalicKEcxtVdMvmcpZh3fWLoPWxklvQjvbhr+Gypu4TnZ6X+2WKvNsuoAoV5ZBm
rrX8naeEmAWqlgO8Xn+H02SPA18mqvHJKemaeh50633DB0fYPWFjEABTp6lwW1oh
6yPYh8ObWxMppTsZAumDn2me5aTbY8JbB9662+wQY1fRYhjKM9wbiXfprXkQwVYr
coRPit7jxFmZWnhCKkdKM0/t4YVTZo8qJTWWKj99Y1H9b5qAaE+STla1ma5moQ9H
yOPQuYCemPjAla6XMHWQl8+nfxIwE6eeBoiubS0UnMv5Tt1kvMWQyHnRnCnabkAT
FOZnjrB5ilBP8TiBqWRBit+XIA+RdpNibEbUT+O+edLCMDMmHMobWIBv5tyvN/aG
PbhLgra3+G+5HS+s8z+t5Js4VNhTc4sDAYAmP3qkg45aQ1wrDKXPYdHvZjQgO9XW
VB9Qjl6KgD2rJK9OGQUn9LayZU4yqN6Ptj165KRcOMi4GzWTN5DZtIyebIYZSm8k
TJ721LoiOdvxrF9Kf9tfCx6mVa8lwr2CpMWI20d+Mr4aWJOUQnTvdTNnptmHNFo0
Efj6iNtDe0G1buEHF+hyDcHJtnujOHAQ7068o5JU51JTHsmmiiQO1HWxXLN+VsWj
LMjzGSmHOZm1MvVcurKrKP4jQtxsGHTtwWf2/4E3yIrK751uQvPN2FSz+oD3mM2S
0BNd7OQjHWzytZlz1Ct/SMQMQWu2jyoawsO93HI+tgTejVOX/h0xOiYO/nVLIkfs
bJbt1h6eSod+VYFx7orVHgDCcr0VDsDlUHjI+7hW2XE5x2z1Sa2Nukdwuq/dRjOQ
pdIJmJvKgH4KD0+weOOQftUGoe/0Z3oiKvUXrbulSd3N1iRFVY2tS/t7inOg3tNw
DdNlt/jcZB3ok82oidMYQyxWS+4zFtg+2R+x/izVzqLcF+1Okhde5x0cHdDubiLN
KPVJv1BvbzB2JVlZdKI5WPoqezpXgc/w6VMiEZCxANR4SmlB8R+a56DKDZEMremW
ZqLGELLkXctMNpAUgSQ11CI6d9lD+iorGc+2qgCqOVHT89eqVoACJga+GFqARYQK
xj5mKpmlVUiBYTfhDakqRQq/S1zEzBpBe5nu7tCNbxMVw4RjNnt2Uh3fR6x/hbb6
p3wBv3b5EgCqhA0jI1n/h7tYXqPXl3QbH80MFkoZ94AjmD4JE9VmbgutrU3mhNAN
fPzbLGXY3Hjbe12iJDcTDp8jL4MyiOi35FX4cC3wn9dKC2i7474mW3QxU5f/VWJi
WwnVOmAootfvq5aKdLAGE4mRnh+Ec4YWHW1AaOrAcHoSJoLm9hfI2sPKjRmrivcn
vHeLcxA/9yvMwfhOS1Xx77VcHEx5apat4jGpJmX7zQoOt0s4RFnjbU9sQc2F0IUs
rNkp8tI541nueqvFaAa9bjxqvjj6VS6frIJPH/KNIlhMucvmeNLa+rg83K20JiND
yBef3Xg5L1ixyN3VwrzMEDazQFLVH4qb5fxgs/FH26She2rgrT75bKfryrj0RiVT
tpHr33PDnOb9PUSoDLInsd+mHU7xp2rUTPafdJgAHI6+oSAt82OTPOh031qDJGNf
Hy4zqcAxY7j+R8kqfIgDvIu5WmLyFSxth5zXG9xFYaMQk+EfPinNhtn8W8JRAquk
4agZE4KU0ovF/Xy1/yEfj96mKXb5QYhBn1d5PChm4lQrVpjKnKFwCwMPfn0sGoMH
TNYgUvtD2wWWnxAxbYBkuR89bcAL2eFCUaicZh2HY1g76zuD2GpgMXHnCwos9WnA
ZhGklz/LE0gAKnAPEdM9CdBrQ0OX4hNfJtC4GV2bVhaxpgnzXl6KsjMlozslLR9Y
C/nRNPOfe07ilmMP3ewzPGBl2mu3HmnZirGXuFbO2BIa133q9huPl53ni7SbUAF/
v+OrACl5+Y8dBkgj7WBuDhVcngfm+AI801/pCNMhCtkGO27HIEVXICj0uf0nm97Q
/Pd6cxN7ASZUS2bFKBq5p7jOJx5bFtBIqYC8kYdQAVtDOvAbMcjwGgkuHaGUVeOg
CaPb17kiFETSDTarWjtSCF3rTdHBYM6NmgZvp3KET59rdqappkjB8/hI+6ONC8r4
WWX/sQqekU2KIiS4BHr88ifbshtS0tuSkMrC0opmwovVpGqNGLaPM9KxpIUnSc4T
hf2leRjiH4T4WZbctvcknTlCryiqX8VE/c30/mrSWTq4619d1j866f4S5534LD2V
a3+TEeBfeg8zMrDt1VGbPGrOr56xrKWTJXOl+4iwpbFu8lKzBuo5+SyS8v9WCvGL
Jt1PCN2bvQOpEaxqwkMginlDIk2JurAaQMwT7jnNCZYg72LCGKJSOe+wi5UuSf3P
M3d6YXgNj4S3o9hi6wopWaqsoIrsoFuj4y3t3AyygAEy4QLf2swWSGCVXqIDbmWK
yrOSjiAmC6BHE7+LNCjwAF/Q2nMOsu9wbwBVlWXe51ia4amdWKUdupfj8icdotmz
hEjcMG04VefA8xoIGDK86RaFTTMHmSID0JS9rilN2llE9b7Vm2jmBrjjtS2hlE65
yQbxLjckU2fRqs/06/VlU0+w/KuoXhdg0CGYJQarTeoszwAhX54YynFKmuuvyMSE
idgVA71nOtqjP0xsJH3ZbV0iyyz3Gmy+i1oc0c6FrKvv/E+yDdGpp6e99bLsa8Lo
yfURGgASJxX64TTUEECWI/jZDCz6LJ4FGB1mCqywT+e9YDbca7Jb4cKiSKD0n+Te
opTD5rr78kjxx7E0E5/xAcnId8gUtX13kC+9Lx2shv6GPb78JBouyZMKLObWrEIV
p5HZG7iTQfYDO422v3OxNVvDLxSp6vOzCpHm4QFcrsW8N5PyJnaYW/+k7N9gFgI2
WlMjnrHHqhuLiYNAW3EHt7nlvx0sLkqPkzyvfFj7ULfn8u1u0EuADMnrhZmLvUSr
r+PNQmSwpWJbxabMBj+2ZDe3Qf/c7EsGpE1fQEcGw6i674X8nHVn/VTydmTOVExt
F1DWBZ64SjE8lavbHQQlx9IqRCz/q9GNQR/yS2yNtB/eT/Bj0O6uWRTD6AbJXZlr
V3eLFTuKw0gn5V3t/LBvMRQLJRbeiMJpmOjdm58iD/Jo3LjmBt2QW1WeQUVpkAVT
xzxSMiGgdkSbWLt4OwGmz9oEAjCSSXyeHrONxGGW2noW7S2JQGaWP45MdAuXucOm
RsdTMeAmz7U7YrhB7jT2p5zpucrAIkXhx7FvAqf1YPiUnkt4uJAzf0Ho+4N1oTnJ
XIhl0HTjwcMeMgchwxAr3IKUm4Sar+/xWR77UY+aye4d2rS5tYqijWeVC0RbyUjb
UjuCcqgB8ksBG7K2o+xi6H4ROMjHT2h15mFWJmY43IoGUddG2OnAehC0P7Ig+BSe
S1ZLdq0X/YzHLFabPFIfAnfJooGKM9c82Hvgl5DSm11FDKZtTYU16I+7cOenJjA7
H1JfPLvUfF4B5PQz5FAixp0JXm+wSxerOMpgYWZ3s/tgVD1INqhOIkhi+XO7ip1f
jiSVcM2qSedxyJazinB/Jrb/xYHwNArh3gbcsQHeL6EHLuSJs439KuGbTGmzJ26H
QzmDxD4IA0LZPKL6iUfD97ysRp1KmyIrvBK1TIE7ma/fb62iy1q5fUNLtK0pYrG+
8JFj/4B4up+QDfGjBTRQE2hiuebt1AzevIR0t/3uTOpTpg6TQeSQLAwZzA8ZYRsw
iNqh2tqRKjtO8vM9vly15NHe76QvhG/wj6H5NNd2EHRckfXHV5G2QgCpBd2aCQIl
u1PNBphSCZgghSuEOFEpylF3McwJ120hY8z6punBisOWM/KbjQpDcRrG9RV4tlHt
gIMxhQPwAn9QFUN9QkrIUpfVRvSz0zKuzc5WrajaHn56CZj/qomMIQy2yvPSE6/+
Xu0AFN47Igk02SF0SFsFHS5IoXBiHsNWERdB/on9mP5z8woa5kAZYbdcQbANv+FF
7ayABngG+VgDfNec9cLtFpB+s0g14oMaXMstVT3kLI7NGrb9dlMi7Cpd7NWJLcv9
n+Nlx2ILnk5tzLnw6PhJlUe1rKheEtVXE7BpfvzloBV0QwvQeNGO2WG5lUWYTT6I
U2fb29qKIORuWw0uO327WpCCaQhX5tzwcODRV/lYLUMOUYtlgmBHyZ6NKkLg51AT
GbUSCKoqcjd4PUVkjHdGTngm1FP9FFmVXdmDoE6j7uYe5y/jr0kvMnZDsLNKXmA6
c7ZrXnuULgICj9Mhj9XLGvAXbwcIvDC1d6cIU0miQoIJJ1kV/+bFOdFZINSMU8SZ
DU1X2INFd6t7sQUsDFJKbA3Z+9QzIW39rrzYWvxaPEWTCuo+yYoIg940RYAc5US/
189XNVAUyxG+bD2xcV50C4mSONmHv4tc9+GskTiNfTBJhuYyFxTyJwpQ073nOcIo
e17SFCLH/89tWHBf3sHGNsupHOs4Sjg8LU0Hutmg6cFFbi9gAA8g/9MQdeqQmj6M
ZwPaGi4L0sHC95sBeItf90HOjYUD776pTseCZPoPq1Kkff8tJo0vP6vZTLaYyUBC
EuK6aavo9MRmddk81EcCjV7mcwQvtdyFVxdzKQc4KUqp7dKNfV5kiTlAT4JYvdg0
mXapFbxxTXp7D+FsEs7f/IT6lyGmAYQp761fGA87HhVhMsyI3XHC7UtXu2lf93j2
Ie7ZrI3nEopYJc83EV6VYNfBPbfo1idJWY2edUOTI31ksbsuJulYxiOtVyqiwIGp
HIoCYUjNzGbCAxJPYSjATU/aofYuEKREuF9c6qvk62BXBmO/c4186tIXtAxG6iBE
9HdhJQi8V9QanGLQs4OcY4ZMkR0guNVOrGqek6vL4uXLMe4+BRVTni/1hcHtjju8
4JV7+RGZbmF+fbUX7ilTaqW50MlxYC9Qdh55ndMgQQTAyOzpMsVNie3ePCojcCJS
yK72uT4lpvvgkoPI36ynWzenbfizoLOq2GfX4iuEiMnv6OIkem214eZdyReLwSRE
l3+jeIK1oln4yTjs56iGzumw6/tQTbIiUArAFUiQ+nwljB8dh75dJQKB1nL4gUmr
BbJryMvcTi3BuNgocCvoW1hpgkJAynL3oSVCa5SggQFGUhhwAqpqfxpKpBIDp5Qi
9etGAUpfIrh0zl+OyE3AmZyKc3e4cet66IPN7i2qLUBFst5YnV7ijVkNcn4wQDHi
1ANYMpUdHj4dw255rYM1YXkQj5XvhXNtSjxQsXUaGD8KT1i4x5+T/1sVNvWs06qv
N71dAh9Blo4iILGrvQfYRgvQS6dS7n12hb72xzklGdZ2PCuqMKqiE1VeLeaia48R
+AxvxCCw2NO6G2KR/jJADQkrfj92eJXhwzlKR31jM5Myt0Gntj1MpHk/6GiHjbcJ
t5RAtMdkhCBN4Y0qFndguMQinCZLOxCKYSrXiYetG4O7cgvgD3ASJ0P+jA8br05P
xPrHmPzzymVqAKFdSV7TFl99OMO1apOa4qa7+xM7DXBMe8zPmilMBVYh6R1dLFnN
bJbXQbdqwRK1oKk8u/uM7DEoYUwAjbVYVteFZm+9uUjH0s2B+OofCN/u3PMHLiNA
5ZrhV7bH+ScnXhRzqzvvQBLYjPrjeMhSiErXKhZnd860uaaDL0ZLN2NZHlCWdugJ
REZkrBLLSr6ehBGXrLoaBmYZFeJXwTevXuW+7ieE1Pt4D1RAmtFdnvR2jliar3V2
trs4tZxr/KIoJPStZk/3GTg+UTuQMAtn4fUTxdPk2Ycq0z0U6cT5y8F+prGPISDB
gjz7e2hEC6lKAPHRR5cn8L818Ik8q7N/GDl7gGnCGnNLNnmYV8DzV9rS5wY2ZEkD
PGz65898obXjUBXUdae7ei5/ykc8ih8jErX49AyPJelqs3g8gFjl5gO1ySUXzteJ
tWBEsc+NBXGwJR5OynNynxTh/JAj3cbAe2qgexRXjxgk3qu5mIFeK/Sysdv63ETl
1IR4sPW4FXshWeOC0SOPoY6icMXc/hX/tsC3afoXrDrDNA2CNcLdnbe6tGx4mVr5
1heu8gYa2TXRk/FrpTyk/0IwQTaBtf9OvQsXQV5EIAouQJoxZbkNw/SGh+DF1OhS
x24VI4nx53Efqp6PCL08qU3q8vgITo304wom+EIAw7WsS5I+r02wWDU56AiZ5Tqn
3VstM6EXGUCclOABithGamKWKpkGADgaf9laaCpixQaB8+CeLUGuvLdxSh+/Ihnf
nD/XP/i/HVRT1z+lcZrLCuPZz7/MN+3mlwr5wVOXoKtK/1RtDBGcSqhlWxaJecLG
BlegxQmEaMYO6akfRhWJApVBY97sE9rONGgS2xtapuRkhV091RcDJdLffhkVAwg1
mRGcYfBPC6zgwsbrdy5HKBo4fN7b+Lg+KMxtfDQUhUc4GcbREMLdzCOsPoTCUNlN
kG62hWCe3rB5gboFKsrYnJmwJCd1iQ156vHw3HnVNY+EbvFj8RgGtdMp9PHWJwg7
qyQAMErkpDhurE0PU8YXkhRZuY+aghW4hSDKasY1422h4TiPflyvBY6dy0JS1Ovv
tIRoyPPpRXCAoawovuQb2+/cIVFexoYkq0Z0FbuLyA9kPm7z47vkVlh/5vhy8uKr
Ic2bKebRNuCrF5seRmGFVw/4O5jpBzXa1888jKQJHieMiPR4FDNcwl3tMoMebBSb
k99T0VlBEszU4S/EalqUitU0hWUi+NLwJfwCDP3vXYhfIkV32aBfgVHCaz/wsa/g
joDsOZJvbri8rOQrtkOauwJ8Mzb8ogcP/Iu6o/yAxaQjMVIkbWOo/WtXkxivBdj8
3Cq+eZc/36TyUkT7ADtyTpPcCZ6PtjBrcfp3SaZfpHDnNzjwKvqhhtFHr5bUmQTC
HqxevbhTVE1eR+lW4fTAs62RxktIj0SafGLytmjKrVRO506YpR1c3oKNF7cC5MmL
DqY8PV4hsUYVzGXrYy2otNViUlKwQh8Tpl+ntBG44SdgHavhQj+osALzVmVLpodg
jKyebV2mWBOzY6VHd0wURZCO3qKEJ5/7bTj7xO9BsoyQ0y4dxZUyrtewoEhf+CTe
aZIcQX3ms5LUjqFTPExj399yj6Ovu625YOUJ7wbNOJELaN4PDShXOkvk4JBmAXdf
5XRcUXfNzC6YeVNseyOUrjfgrRqpCCrlPcXZIrJE0KHAPhbMOSttJNQ8s+HYuEzD
Wp3cOTQSEAFzcjvaNpVNGnMRuJ0+SLRBjlf/U3SYZGs6lpjD7mkA2Oru6Eu2VB1f
f98VKDqgTgGwZ8WObMA/KGAP3pUc7Mb/ITMHO/8idsAD0L4+2OWy02NUSTBkk8ur
eDqgaCASq3rYBJcGBXA3tk8bs6LCD7mSjHdMz0s04QIktG8V/WtTU2pdNpp4bBxh
hhDN0KMpxMOAGxB0ICxOiaaDzFLGIgkpj6DHL6bkZaCLN6D2a8NkKV4hgaLhYNXO
Fw17lJJXudEDDV/n8cTeItDsSzy0eiqigCyNEOeeF2KRIRXS0nu/zdsg01+yjtui
BbMyU6yhMRATuhF6uS29ZsksNk95IlOxWpddhIVa3KkDA0bafqlF5VRThCe9wNH7
nO+gFYpF7OJ0+eKfpnkBEJ8QPS6HdGzAe7NDIKF8I5xtT///cmWb9WWsjrK4NmSP
UgDI1leNDh5tmM8ujbyO5zNJmkUbcOU5DuvyqGYarRQjokjKP550ocvBQi5B/uZw
EuWG/9FQT37SzEAUN2JpYmvL4OEkXWX1O0WFaOqJAyh2brZHH8YYkL9qIf5Ga8c7
txEOFX+HC44r5T6wCZsBMozXhiXQrbJWoAcIaYFQ6b1xatVFgUjov2Sn0sbSjAoL
2gTukPMqszzS+ZDWHW7P4ETYNXEtvHAc9AoT1c3XSlYcZ1eJzAHEH16fTk8NmAEY
5ceiahMPH5WrtxUY71/2Aij3vBDTc+q+lAFzNLTj1EihiJhEXResNW1NqQgZ6bmP
/DTaRE6qe/4F5JA4rLSdQgNNQmywNSyXQ8hx27Bkg4yLykgnfdJEyjQdx6sKnPaX
eGjgHvahQhsTgwQpAMryhmM1sTyLI7KkpSlzmb/hMXYoI+KbUy9doKRz+f2iNyzI
3pErioz5nYOWjzCetP7prZUXurqZj59Lr3IGB4N0bjr8Q26TjsRybYIs9Z+GpvBM
oHckZeaQpYRi7BEc9HBXISPwSJislEPOOYHpxBYEtIt31wRTe7hyqwQXmt8CEzNk
bv6zElirbZMNvc9iehVv0lzTTJKwn82Cb23FGdJBqBgWmgvgL8VyX/Ga10nxKT9h
CjM9CEJ4vrkhnCBYDbMn5/erzv1qhLXzBui+QYfjhJdSYvvbPGt+JD+IWmSKeO2E
2v1NqobvD8WWWepv2dHGdJt2hbgYPnMgexzt5Ek5bqw+dDKNHhJ2twbFg99JcuJ6
kb8df5iCefdR3objNlomeTL16dHqtMkU3beMbvOmsGMnxrROSxQv6lN1HI8tA9nN
47f5Qktny6m14Z4lktvGmNYHf/Tcj5xK6vOb4JM0HX72PpzDt+jXssAM1HyvmX9s
n0XQHaROVARSPZDzB5Z350wjmiFA1OUKwmYS7GYLuuf5nyAW+BHRe8EyZIaq8gGy
NtC6tdYG8j/JSqNGsS/VgBgVY+G/44pQnPulPAufw4/EejpRqL/gFB1hSH2s6h3n
t2xn6zB4r1x7IG3RN3448Hsr9bF3FUcsCLZJMoUndiqFc3B1dL0dIROLFX7emjYZ
sd/HgDAtIu34qFI228fbnwvFLUVEyCwBSJubu6ltR4t7H+oJbQ4y0vzktwbXZP4T
hywfmMiSKB6pc7MoT8uyJ7dtkibmrgLrH9MHrcrIhgg09jwRctNJeO5RS78LNgTg
fAJ6Z9QO5IM27PfMadLmMD5HznvF2LNGAaoj/I+lm62rh+Boo4R7i7yISYz71Bnj
+RisrNULHPfcBcF3zvMZtDFFu4KWKCaMq43speEMb/vmqc1L4BlK1QNRk7vRwSq0
a+O+YWMVBps8SY+m8ITiqivAPrUbLWgFx3bXp5XZnOKTEkYYk3PUAyIM4qVnM3m1
y27jXvoj8kjQncKjidi1DufjMVajp0AJts+yB5qaxCKqhIXyGHfzN1WvxeFBPhYQ
vXHKjMZ+BIPrcEK47Eik/qCDIaYIMccszwguXXDEJqqvKHWt6uv6FgJhMxHUmZHc
v6bseADhgkePah09BqAOH87aS/zUvZF/8fIUHw/qA06uIU112mh7zC5+UjgVUAi+
sTDE96YeiFdsIwpoWqnTtdoqxqlGyMWEJOQ4jpf4qHXlur1VRIdBCXwgQAUrHnnm
33CJpFAROuobjG7mUBuCpsB/zMrTdUkL4A/QSIFkQUf2OvHbjqnZpQGarQA2zzCe
I2ZIsPm8017rPWMP0Y6YRpvynkXG7IHdKxiBS7S7WpSWcLKub94yqFg7PKsZ8VdS
1Bw14ppm0HQhX9LVd0oD3ifBACh8DTRO1qrfINwXaK4yCcH2xpesiN7gcshRxBsg
K4ExulxqPxbxOZlC7mZIsBmyInIKSar13HqFZX13c2Z3BJk9Btf+PFwy2CT2Epgx
pHisDsazeEukLjAZBSw6huUCOEkG0NyzB1rasCbdz2VhAm4zBmBXQiSo+WP2A13L
2qkRLuGBbCbI+aVJ1V6N0uTcZISU0YIuI/fMTpq1Ji54DSRjNCMJFtrgKMvPsO4f
tGHMC/zA8ezkGx8brqczhIsUB3QHGmpz2AC2BcwcmfKbLjK2J5c8j248w6kD/9DA
yyxUa6ECW1mt7oRmTmIzfcfzuhuHNs/m3wKLozBx2VT8PLozACzhU83r8OACJlV1
D1iFB9z6U7M0ibLg8jPD5kmHBPnwlAlz3FcNaicxlYH5ug+BgsepqSzzxoHd/we8
MBSD//LwBpYObXMlNOHw39N4thQSvs+jlAUfYeP1+aFmfTjb58127rE5zowYmSkT
hlDbBBhFIiYy13IlZtzj3Zkl6cRzVfg9zY6qECOgk9qPZiyBfioqQH0nApd4nY01
a+o3NyG40XXyLCZVnNMEl7wyl8oIBOVYswmIxM2yANxB6S8/Gi8LJbKD9Dv79JZc
rEjI3tKJSar4C3r5EXbGddGr9VpM4TR64wi2PZjBCfvCyorIYrJdWCMD0jFidmEE
j6pyGhRPBhlmA8osaXTpxDV4AUF3/WN0j79K9VvPUk7zSEhHvmwzLrv+doI7gWp0
manjjz8AwFx9Q+9lK/tMRy00/S/bFlEBEp9gHgOX2d1upkbe6KgCM2pyW5O9I3Kp
r+FZxfHqz07WZveWsnEeXkXCplfegl8Bh/mE4ToHvzbsqEI4WzeMgGGEDT735ee5
4+aKVMsw0MfcWEs0Mv4aaHkkHREZrP7plEWu5y3JM+6O50BisEvxxQUX25/s9ZaU
cm656XjbRrKTHpG1TSCT2A9r0d3Lx3tIzp8vs8XbyiPjCfiKAnB6Q21LFacRV5O2
DgwSscLEzWYwX+PAvRXufIjxzIeM4ep7Ob6+0Q8lJHBLtI7UYJ6Aw2+W5LYi1hkl
DSudgYpLulU9NARAaYk6XX94Dexwa0G9E6tZaqaJxwMJu3+W8mQM8iK+zTCiVnrm
Pc0lJd2G0Fkhe5RlWmYfb2prGiY/BtZ0jKN4LbnOvs10UkAs5A1nexSQrCgUkmi9
5axXGMpVJvOlaOsGSaf7KZSkZQolNJvUnlVQN3ccG+bqEo2q5p9gfQ4p7O2EXuRx
U+phBsDE25E9Wv0gPoT5BMbUMkBrEru9jb085NpuY2mOuz9Fg9eugIp+fpbi08kK
DGylo/qawKr0LgIwnE4gamrQszPbTB2ImImVP4KZaNUzQTgHyYXdO3gDZybcfFQG
pLakwNgjp5UwAVBH1jmqDxcuv1z6SUyLE/Y3Jg5eonP2+D4noxfqH2ZKwCShzlRH
xf42ukxLJW45Zb9DnAgLrjPbtnIa905/dyyznYyGRjMxQxM5uB4e6Duk2nyg84ec
yJPA8trdrL6EBdyRA+hGKA3FMsfFW2kdLopOYNf4nufqxT422gSX5XFlIvCphcZ+
1wcZBKIPq+0IXocpeWgIl7DmKYMFKqbtZ822J/WNChwlIw8aCw5yCgXVSk1YmzRJ
8TivQj2fHeKtUB3ykLKZwgsdE+ljI0HDF/0oaS5c3m8C/ofdIBwjjXTRxT0eIniB
Ec8S4v0lanj2hwyQk0J7Rgv1tojWMhPJ0qrVNLw6S6gzkpscSkMAFBjqIsrHmcLS
jafEixDTWP/Dt/i7hpc22MlMYow8x0szVvNTeLd7Vk9mcBFT1qYrrCPJv2DBTTIY
/E7IJCC9DRSegqBv6gtHzz4dD/1czfbCOGb943P7BPpXUYWhu5up5daNY0DbJCor
8B1SsKuydqIw+qdJbwt+RFABrcWN+NUQy2jorXUcy0XUl+4CupjzAcdbjQa94qsa
b4MssK/n9x1EtjpQKgUylV7OTQl2J7anl7dO2vZTjyhgwncozlAiPJVxbwTIriSD
Dpm32VfAOTP0qQvovgLS1ELDr1dVSDp832bt07Qe129JTtej/lLbmURaz5v5ApOi
PgN1v11LfQiJIOnrTOZxD0snbbkFE7x9VMlKY71PhuiAnNIz28LV0fg8+qpSmRyT
Q1rym82CKtBreYHLObWZ7l6lmIL9N0brgfujvLh3Fn15u9hkOI94oxz/MhsvmO23
wgaxbuZ/5W/yGuwbautEPUbMzIxyKoe5JNpbNHGK6oSGSRM450rP1k5zrnCA7mCS
5P7bbjmReEgqaHsGrkA4BxK9xJOIk586giAtBHuzWvOppCbUnFBGVrt6REctIdjr
OFyxWHB6+kb2ajuaoAErXYB2uA3bi3eaS0BPFaTs3KylpdRzw+QSkjqFq3m58xLC
4lRj1FuFqU7tcw94wtFaanrDtlJYQjpdrGpJSgWzqK92fMJKafsml7+ldhtrufO7
e9XcSRQIvhUSBt2HBLI7tfRI3Sgb51xIwa+z/t0HOPlCLF7YwbvuOTxSVJyAXENv
OFsZFSHob0Uk7490428cQ0h143uLVKQel2uRHzHHL77Z4W7QKCGo9wje2nN+h3rx
C6SJAww8Fnj5nWF4Qw3wBVRjoR5niwJ9FF8fRpiY+u79BMCks7Cg4gPg8ZRVaKUP
BHnd63vEhdIxZawCMliOoHVB26HdLn57l3T655vrkM5Ssok8AYLNluvSNbjV95yP
2RH8fkf1bXmO/KyLpGA/Ds6YiJ/jki02Qa0m6fcJzYsB9R56V+pRBrhKUUz6Tc71
qBUj2E1e+orZJfXQOC/sAJtcmKInBoG4Wt5k2fYCd68CESqmHKlkz3ED2Zw9ppJ6
UqPvLuYFpKoMuNKZ47ZjLPyotW3wj5EhRgPAGEYFT0mvGnIC2nvXLi+td9wNyEXm
K76SYOPstf62849xRVHSECuDGLZnazSZrg8XmDslojgdZdsvvswZThXT/pqK/xzT
aQDXOroA2yUbPAAaotrVWahIaTJkuX/tMdBr54RZdfjvYjn3KSPJs4RTgaTVy6IR
ycz8geitqqN3/Mr0ABP08jQlYcJWnYr/QusNUA6cNa5gCb2kyYA00nYXeAAqaEU/
5Nz/9xrrF3KLmpIVy//19or07dQx9IGwFsKjsbGrml7O2fJuWHs6yv0Md+Xb06tg
2287odk4eP9kzxZ6MZR2tqjzcKtqZhW9wDj5aLjJe+Qenxn8TUc3d1nxi7wVbjip
tTiNTdAqgvMNYTXSIUtKLqfvH5BRRhfKy6Q0LqKo0wd2lo0KcI6npTpLEpq/3lxK
82sJaDr/fpDgEuYbDg/NEBNBfHEKyDYdDweuGDbLiOfoRlF8koL082HK3oZB/4Ha
ahPoy0Qiyvvjr0l9RhcmFPL4QdqXamWVy5z/ch0J0ifWRteP2FE2v6cmUcbfuIhO
5CglxU0KrhEaHcxy7vi0EzSyndD3zVRSA7ndtnkMvOFMie19cHO81RkuqCUIOpg5
uNRO1DuSwndpQOK33Kl+eyfND78tTPsOX8wJ7tP3iXmVpGu+lhPxRy1XPHm6exqq
SrftPINzkeS7ulX7763iHJsksW3cNe2iEe/LCOVP8253OOIm9y/oNrD1177sJCHk
ixebvehfSP16aHm5avGqGznu0jFoaU6ONonV9I15yeThrErskyVSz/dlDSTE/9s1
hWhilQclKwmY1gXUMcTsXndi2LaWPA3hvSo53IgLHPssSksyZBc0VwG6/JM/1JDh
7bzVwr+7PeGa1KmxQpfcGuV/IjSIaFCnPlk8tY4A6N7j6nV0Nl6tzWzYWHsQAYVV
0mO3RjKMQ8HOvlVHzy1ErKnO+9kzwJ7fZhW6UPsJ7LJYw9BObfWiXQqKKcXpwo+6
bmHrkBYW6MTpvZTYOnWjq9SJnx8BNpXlA+Od51Ebb7Nioq9xQCJLVL2k5b0ryAYy
1br2ZwlP4nsjiPk5KqIq0azjGoShIXsyDRMx2KSOCoCjPA8oa7nQZBVGkHbMkdwr
bO+bRp4jdQhqJTLP6OoHcPpT4pQksOZJbj0iKSxcaWqo1sSHS7kixDx3mvD1q6Fw
Fooqn9w03Ds4AvTQCVd1JgtkFM2/wudUJhkxWWxj2Nsz+gpw7TCU/HtPyqBA+uZz
D7zkqWOoqfsNULnUvpkA9tKVF9DOAy+sRvvF2RWhZIuAV4u2UuQ1bnFyJAf8y3B9
+71AvtHpr4TQSlYhmRu5ckKToAXp7dETkDFx5gU16ZsTnxtj55TqC0hXoqM9a91S
OtSwF85PIFPyZUajy/MbaU4XstbIUZGS/yaVU92cwKl8+j03PSg2Sr1rrO84rnCR
TTX7+OIwg3s0NGJKsxsf6aUDMrfboMWx/iZKaJ9jh/p57P9d0g9s6rW5BxWdTSAO
XImm1ULm6mQ2/EBeqJza2U7ngtnsFUa5TLC2wZ+nOfbHC9QQTBVyWKK1dyThxzmC
yOHFHy5hGXQIBaAtUELBU35z/DFE+ZKNIQil1vSNlxcRsLpkgFfwBCZngNwuiZtM
en3OzBzt0QZRet2Q7ap4zQRQ6IZk/CjbXXoIN56q+ObQ1L122ktnJKVF5r9ih3jN
U6GXZndCk+/yJkKI97DmXjZeOxw6q3LxCxd6el3G6DQBOffYpZ7jb3Igc/AGW8HV
IJrxmEYqeMFhDNiHNLVJuSmRpZYN5PRBOqJbrRRAJSPx4f7jJmzb0xC4rs6guiSW
QtEu5oJ9qy9Z9R3R/hRTego2pU3uLhEp0Wy8Auii/pVBO+K7SY6vdBMqSAZi4oLH
NK3A8DpRL+Xz5NFn00ypE+ItBuFzy9beTzjhu0KFVuQyWijFqdNZrUkH6M1jc0Fa
bcjgosW8Y+2ZId/OdcM/8894oTSUwRhuxSwlVARzZ1ZxLbnbaJ3LF+gfvUuVhnDg
+QnYGzLxzodGkUeaqnlsfyJpalzhosSBLK31GV21W7FFdi0w8xKonJgSe/cd4xQ1
TqXJ5LX23UYa5kPOLsATGSqtxDYB/2LMUNZ6qzRqw06bYnTAqvnRnCGSIFvC1Wqd
4dhWxHkKu8Daeh+E/cQfc3euRfAggVfxuY+PbnishXrHBAy9FRoLbeAspv2vinRv
nwSKZ6OY68DdFGGa4+3aQiK1uxGfmlgTjP8LSFGWwe0sbN7XN0ZVmiqIUvtVKAr5
Q/+vEU+zLQ/o+9zQCIUavU+SHCeR5wSyeHGE+EL7eOnil/RjV2fsKdD90iZEXOpd
UpOqUnp1i5tsJQzibr0jRj/ze/T6eP2EtRYuk//6on05IM1yo+G/nOZ8BYSqG3Lu
EsoJvOOnoVByx1s5W3iEGBEque6uDzQ2fQH5FDp1V+s/ZF4TzB1Es/bM8qlLIN78
qMBTYaCAWkN9hKD+ple/UU51Qv/mhI4zy1MmsqekLYnqi7g3DPcC9P8LIiJpuweC
nhGlp95N9RhnawlNKz447p05caECINzk91nUIvM6+5vE+78uS6zlDNaPsRTowAxy
asHHOK0b5UsjEeNbOzYcF7SDVzcGxFcBcxTRjymyfgqyvyIH7mpZSxGDEbWkb2EK
tzB+cg/Kp5ZByoGmUhC/Ib5cHEJBMorz6KkUL1OADPzWPA3IXWW3n+4glhH6+s8L
LLfeDo/NNZTAiVaWOk/7+gqkKop+EQgSYcbTZuaDtU8H2cOMAcpD/oDx9fR/36ID
2pWa3W0kU2ac7p2XsDWE5vt3IhsuXIWa4trn8+62KR2iHurG0eN0gtLMH4uFVBKc
gFSQo+MAcUs7wfKuzIBbPGdH7vrQ/tXcNBdJjjEBNYB6Nw5acCN5jNJzrbqyAT41
IepIyBhtR0gxd5W1Dm0hfXdw646LY0ULH4m0934wzg+gzvWSID/04N7C4X5hTBYC
cOdBBhbWy0tB2U08tkm2qtJxCxFsMpHwdRX0s25I9FYCu/5Ene0OAUvYcFqmx7na
kXpQWtS3LPx3NtO8AXX2jhA1CLyW6iH43U6xZFHuoNpNKl7rv0PTEN21BhGxXiX6
8LR5Rb09VFEwLZ4ZQgi47h/cMSgsaWLei2lkHXpo9Nuiw0YT4nVsfWrg8yvrfQCt
ejBv9MllV8ULBYVv9L1dEIkDJ70qSUFkSG4ugbJ72compkuGXunN203I4Ru6KGUk
aiD0735zFCjYug84sTLWUI5JdLjPkX5vRyj/OtYhbrmG9pFE7K3KkyNOGVIV22Ua
icZ/IAvET7GM3KOdroCxOPwTDeUCIzkvHld0ZziDAvoTmXHWdpiDsxu5vZB1VvQL
DKar2EIPDHU0m42gdYrSPV7ahJp5Iz1NtRjEweLBuw3HbekIey30Ei95gX8UD9LZ
vZ9LNDRkOxTnbFqFlilaymM0fRJkLWIXf97ioQgX5NGTO0RASdkwrlrS96+QL6dz
rsuB3TJNCvEjJlfR5Y13huAMf4jFqq4LjOwJTW8ooejdWU2WP+ETiuRhhoYltgvw
S4MPL38TYw61ZEUbNF/hlPW+JZzmyqkrJ4XEzynGEE+8MQJUUv7LLJRj6g6kkxTD
khqq4oLrEUKvQc/lpy/3d3og/F6AO6ZRI40JvreHeUOkDghUn8LZTzoQPnYpzQnr
bPSRKjeX4q76z7yEal+jr9EbilGw10ik4Rd5NXv3LxmzqrL+n/bnVivziOa8cX4M
KtEiSKaja1QG8WWnHmGfdf5AfBmqONCRQn8hRmh2G9qngke876IOR4smGqJBDrfs
EenLD/izhrKxhYnBZ+HjBzy1avDza7GOAbUaU+N8dIgcAFGafWxfGXVQpXklBkxB
y4lrlxGM1inbyBiWEMRBzK/3KUEO7hgowlFS+P4DTGMaDvZdEPc5mQv0w1k6WCLO
THodY9q54nJRCI/RUUWlJPsHa604UVNUrvCH1oKVZnHdpZW3hqUBv1WANgvwTGa0
t36DGwvkC+Ril6v7my/QrNoyGkIJ9gRBPSzuhDPCShhbWaUphxwT6vyMVrqgX0Lx
bzDy4aIfSVhI09gvD8lNu72zv8d0Es4jcYLUjEv9gAQ5OisZN8oUenyAQWxHMhS6
ty7DjRM99WEzd7MW3VZ50sCETwRn261KTdFWEhn7v/+P+Aq8q5ZMY1vqShRj5YKW
Zt4e4+/TA5L6a+dVu7/uiehigePEW3svwIWvEn/+xUaNhHd1NJCfSjotiOzbD2za
Kj5IZD6Ac9hNGCwy5Mj8jdou8Cde/Y3CnxZT/GD0v4KkggWFaAsGGULP+gpKS6o0
u9gkRiGMbRTAO2iddncY5HaTC3vC4aX96iSeGz3RHSpB/grXXqXbbVulECssW16S
1iloJUv7WY72Qp+uXR8FED0Wl2hL2ahPLTyKjiErk2FY2LAKcu7MCeWjlVzbQwPr
Rg/rKOXtXtsT4ps/iZnCTdeJHcmbTqUwjuX4Y3hVQJ7oKQVsbGIPhmRKIV4AtAdB
hmtc/zX03rQEYyXfPoyioDTH+G+FAhlPL/4hGwIM0gDqZq06iJgMUvmyoqMZG+UR
bdMOLSEUXrllPrlVVxSwMwdGGCG8lTnk3dOaz5WwssHMTml/Zy6RRd0CrKB4a32v
eCrBdokNgMfdXeh/LThoO/vh5EB8FhB+vIEOp+R/G+iAVijgExFDRmDvv/mAznSX
l8VInmMOTEFrlXBuQNnJ9yWm9/BESiZCZk6dXfv0rpWsQsz77yfyz9hy+odoF1Qs
W1CeiIDGQimX0x59RK0Tr68KBimoBBNQBFG5k79kHXwGcNZ2eRyriMgRkSfhQxoO
DmO12CBZNT7OsRX2BjTtLl8kIEnHlqkXO8hn1uJYJrHYv0kl2SVyoRI0yPreGQ3J
yOArUPzCqKH97aJKXBhA4UojvmPwrye1n6nORbDmA1SRJ8XuzEAtBtsSzSOMaq25
A+EQO55bTXYsl2PUM1KXyrDIaIkJmjnq8P5QR7Ve6yP/JGCIihnVWZiaHLeWxvra
vC+/uRE/20HOJPGNj8U3QUeGUn/yjHg+di2B/CQZ0o7TthPJNa2PsO22AQpwg7sV
oi6pV1eLwbuTuSiV9BDyjHG3h1yeT1pvW5L4HPFJClBV15UWoX3dA1zfy8Reigkc
jv/VTCDckF3Dj+9/hfT6kldIlWD5xbhhlsXpWjTZq+t/oTGiaZQA368St5qBZCzl
kUwuLJiEIiaxU/Cp9Mq21hSumvLYYEgdNxMkg72Wf+V8tIcwfzmZQLZk7OEyEcQd
eEW5aTM+aZRfWjoyOLK9CjiDmk/DOVISONVrFoNPUNLlUWVQczLw5TchBtwdCIaw
2cJjL6o7dDzxbdl+rk05sBUIYn5585vDMngXm6sXFcOfMuF8jnpahJtYZ08F1le8
D/Yw2sC+3PoKuGxPydTZKrZR8MrJIbCJDqcJPHyyZaPeq+WYKjgE3wZ26TPkDeYx
Ht+JcwlRq6Cjjw+pWqqxpU+lDlVCzgKBLvuYC+Bg55zW08uKv5VoKNn4o7DnoSM0
EAoQ7RNhuPt0IgQa55yhYzZVHU8qCWf/Rf6NSA+29Wb4EhGfwn5B5rtseLHP2Mr0
CxHFTudynnFW2hXYq4D//TL6xCMwjEhnlIYkJB+01tBlgazSQjTJ9oTbZt0g1mA5
HlK7tFZwk9V98C0BNLa90zW9ytuPUJO+SJXWIL7HadxIdKpShtzzxEWajnHlvb3W
WLuF8u1Y3QwMrnFrV0mBPBDDwRJ0IlMCRVxhiPTmZfP+JfZqNc+vy3ilv/Y5w0ZQ
wAhPEksfNge9YkFBplyKf1REW7XlQBvX7eTWjhBME3/tEl9taZNyLNN8ayT3Jdb2
uEbFqxWfrFbufKRDH0zJUWoGXhzGhVpBJAFotzfMFm+VIGu6q3BQpZwIL6HFFoBA
RcJX0J4JPfXXNOqQEPg/jX3q2JXus6KBgjNEV/UI8FunuVr7XNzqAPqQezOvh+6X
1hfxsRrYNMOiKXLaiyrXg/cq3D+ZSnQDG21+kR0njOJ0mNEN/DGTWWzOii9qF+I5
wOcwt5dXsNG6ND0tBQJjcmlOcd2KHwMrHSBLOQyxHPFAv0BPqFs+4+GgH603i/W+
MkAbWWyQWQ40l3THkIjZNfJGZ3SOCcdLu8oLVXZOqsWEj8k3v9Hq2OmVEI7W+drW
Wy+9jBE6H+rCqJIxAMKLH/b1LYyG64hMQLQ4bG9NxlK3fg+SEeGkCnUpkr74pec3
FsexYsJ/OKJ/h9mh37nICVrba5Ifwoc9r2sxWZfpaMehjq5iTlC9zmz/yDRprmvw
M36jFeAQgGvtW+xRDZJW8cQ42XAvthWqaMcmcfSWnPjgugOD2WX2G/C6ef4qdaVr
7pG5Y0M5sppDCjUZ5UqDA5Qj6LIIs+rGsY0PK3To/n6QrH4LzRz0VCO2pzQfNsQP
uiYi9gVteP3QdigPQ3HKCT7jD1lfTGnwBhR+v2aX9VB4hT4VbtYKk1kzIkB1LXuT
cWFNE0jTf8YUDDQLVwKtvF5fCRPUSZ6YVFpyxAUeA0o+FK50uNQK9rXhQoilgvcD
oYbqo2kGMDY+yedzJdpTXeUgX59kOfqzrcjLKP8PQYk5ai/1cD6ZiU/qWJdEiL20
MZygr9kaaUqpNCNSMxUTb/9GYH/LL58I5skUZjn4wy2AD8TYepvaxiTzy744OePX
1mywvnsi9MvhZg+e17WpntepYXx3IaRnCTs+3XDdi1oKL4YUIB/AAGNmn8ECcASK
D+S4O2I4mnnYmEW7mu/VD5MeCQyOruEJD8G7sJNi7MkGK19bnqu2RKXudXwz1biI
VHNRv+dLV+c2RRzMlWetPROXeCQPgO08I8AZM9fZC9mAs208KLr7GknDOCusNf6F
VM1t8fs1d3DNTYAP8Vg/djjOHFZcN9q9UrduV6KhuXqD1GVM4C1bq4h/SzXHBqh/
GtYzH0kGRPepXRTBYsK3LEpIdBMAe5/svtffqXVFY7hhaVU+Cn7C6nnFpFXMDC6r
oG1VCWJ6Tjdi2tZAkWxVrOcvI4IrEHgOzVa2diJmXE/rJIowlKE47daNRA3McoV8
RTlrFdFelUUyCJIuSWAYexitnDQdvGS6K9X8DA/brZbeIlJbsIRwaAiOXRimcFCp
IRt5NOBmwNxxWlZNKxuWvwjdgYXDW6UzYZoQ+NuvnSwbUgsloN9aHysSnfcj7XvO
LWMbCdLQP0/YDkKQ/9tAtKPGx92uiN20S1x9MPXniA0k1zoVMtDIgYMPKkymXrWO
iJTHOtgIO8j/nVVumSc+tgiTWTl/I+burQ5G35Arqs+mcmnKl13vx2Q/ak0zkjvv
AMUvdij29qV5EfVzysFK673Ljfzht1DhNGlg78VPwCH5p07uJ4P0jjjwhasW3hNx
LK2TK+Px9V3wTEWuq0+eeyuaQDBHu/6n3YW3oTIXtehE92+r6l4Hb22daJ6d41JN
J1co0oWpXKKdsKEquLfFgyT5PcRyyn2z5liT9kdLgcXxecyRYNKvmFlAEP1RTawH
f7mwqY49LFDMG56rLzC91Ry7Jxbpvwjg+FhvtRHZfBmlg6qTHYpPkgeKuGV80/KD
2FFJs+5y8H+F7nwgz6MGq3aFzci58XyFwXUitKQpXtwkFzZEfsocq/vobbKNohNV
lxt7GMdCQibf8+Nf5BeO2i4fLG1pmDDgXUFw9v/jTK+pQRCj1WbFKbV13mVWmC40
nNWLtL02pp/e04gMXjRjpWlr1I4qz28lzARRcKmDvQBb+tcn7xVN/aWDC+V7P7aR
bGbaiLGCTxkgfDuBMG/Nud8iG9cu933vvvSQU2WkRHlCHW3IhHEVvs47AkhXHMDn
gmMLvCLcedpO0OGTVNtsS7rye9wzn6MlZAjZ8l1BHQH2+lDECIeb5kyhGzur9quD
aVr3Oz2X6mcdBs7ZgVbXFTNh8rxLm547CLydSZnektFvis3NSOhFfMuD4I4CVh6s
byuu9MW9tmvLOj50UNm/aa36BmFenBX9JjdGu5ajcfpWJpVhI4ZM64M+7sAxVhx5
+4xZU6japD4UurKHcZdKpbMFGBBvxy0PgLZqoWRzZEGVvQh/Mm+QOBaVXlzojv7e
RakHHZEtHw/u2hpTbKCi9NgXXNvfhkdtwLdTsYHJTVNri3uwckZMzth288r34Am/
pJ1oCHL3Zq3avqv1khW0HK7x7plv/EBnG9EZlp09BO5HJuCt/Gnh3yy4e3xB1PB8
Ybtcd+mUNgjYpeyxyNxA9sOzUeTnJm84B4XXrpovc1tsclCJwhPjEzmw7tXdAk1D
me5VNlEViD0UIGS+tCYLLSkb2fHttk/DEjfQ5JfWJumauObw+vpyJrfYk6PYe8m2
wRoeCB+yU7PMjs2vWg0LRBvpz0o0a7qBcakyp0OCFoPcejvuABGIdFmUIPTftpa3
shCQjb2rSPFOvd9/JvSyfgQsAJsn0t1wkUqgwZD9L+Eoc2SQGqx2swM7KZB57DUq
pfogS6kb6dZ1x5lec75T0zjIMmDbzFuygsh5pEcz94so0VZNYr9/Q1S5eUvOTcKJ
fOhRo/qRS9A/x7ocPi8KQ2jxydAOfXNk8pBsf5cl3gXpGduEABeUnUumqtoJDECQ
ALHWqZlmMLAVqPlduHYQWJojNI0ceO+kU3T4BuOZbFIFTUl/FdR/gqiKeEJWcSdx
9k41kxOGOzhAYOxNq+2S9xZaVdSvcadMh1cYa/tDlSBtPmjPGZ+dtojMgZseLfpf
yAKpjFmq5cuI48jk/NAZARLBgVlGqauctiEq91SucO2yQEMYqrbXcJTl/YOzmv01
vwByKAWFHW7LDWrXyKQVKt36L+7zn0iUmq2Z+M9H28/+CLwtG6+iCa0P2B0POpxs
k3ZllDWL4d8rtjf5vk+6mHPACQl6TYXZ30m1V3x5fEGhXvr+zqQevGQbMICnNdtK
7tfiS3udQUDu5LJ31J+iMgo3UmEN810CTwRPsEHW67wJLLviK/9tQJp4B7m5A7KX
IhoyDGWytal518/k9fqpABLmkNCjAIfPvfPaJIxpoOcU+b8KI7mwnXEAOp4Rc3TQ
t5c9UaLp4wriIficL/5tuZ4EQ4BTOV7epWFckv7JMnRqPScQIOiK3Wq1OJMSbzeQ
vxLwcZQQbfm+sSJ070lhmSeQ0ZIJA2FfV5LOhvMcDHxzra6PKAfNl8w0qWQjEALd
7gCjWFaM6htdFiMjESKO8A4aBjfhAb4q6gJmNPTlTpHxhlLRnuzre0oy2kByXwvh
5rzHjMJ2TSgSxaqiZjfujw84NayMayyxZB4RQQrX1nstoE5iJCW94y5NiOP/TJx3
7hIvUk7SjL5X4pPGnZmKdw1ShnUH6YTV7Mr9GKHPF4wfbUTSc5TjKuvjIokSknwo
Ypc8JePaYmV7Fm7NE+GT7ixArJ3roX43zoplfuCyxORWmgak9nID15zxkEbB5RtI
Qv1d3KUmvrw0DV60cE/jP9HWYO3HudV73zfSrN3AtUocRPclf1y7rZWY88zh7Lx6
BBA2EzrRYpz/qFCgIYrN60DXDx+Ph1qrlAMQT8ud6W8IaxzPDoTDvjqRp4ieCCYu
Iud3HgFKQrBQ1io93nHN9zsVb6FGQXUVLoZjxDiziYb1M05zB66gRae3uHoc7twB
bJ78x+BNneN8evx5sh6TSvO+DJ3QH8Ht1+h2aIfjCMCff6WIV6Xt7JqF5NY+v/5s
iYiOe24tuWT+BMCFtLq8a+EFTNZJJE8XFwdsjt3qBt0wcVE284lDVvpRS+Ja95Hp
22KXuJRNe0ftU3VnG5F62BUdubin77ALJqoX18AxFsRPy44uh3HveyjnfLSHYCcC
lK7Kdv6Jt40hezXcdB7o0ngsdhl4OpRM1FoW2ng1ryJ4tQnWt+2P2ssuOxrfP7Tj
nr9+9JRULJMcKmNpus/ez1L/qNdnC/xpXQocyMLMcqZFyxVEdyqiyfHY/uCx6NEC
1rHNgw5dkRloungzr3deyfLS+QxHKb5z+DV0jkdlh1aAerM/YkzUuIRiKrrVTfMV
chnpEjLYCM33LICQNLJ+Ptz237Tn3Dx33dYwAcP7UYRhDUh7asW4yOiQHlmD0klZ
qNiB9/qpa7yauO7a9/waK90QGAky0gRRKqwUHwilYFoosLMoglpC8VTjj77K714Z
uU+en5dO46pnLBBisFaa+LCLU3S3xt/517+QAoKbQlvEqiASnMkyIxex5js7HaFW
gV57V61TGwN6lyPuPjKUjWxYyIW1VEXwd2lYx0i4NlaaG2ZVG1dDDgrJtULqHqUZ
YKF4jAIcjfJuS4BSyVoy9zOmKmSc+c3M3c0ssWPNwbhsJv/TXAupe+qbAr2Njbi/
4FkFX6xSqJNIg6zy08CGMeI2rBeFSYQ0UfsrhClz5aKZxo2hU5uShO6tTdG+ve7i
Es5uzl6An6dxlS+cqQEncO3m6GNXu5Ve6iKyiFYxHVfAM/z7LpVLybM0X5d4sWwr
XUtocaFaxgplrvOi1eTTqvuzKI4wiVnfvi1gAJzL5Bb1LVT5zEi7qASXwJBuoeIW
OYhaBph8FFsWAkQa5TTYqb4+CasXLnQm3upzKBe7owl9rCrm+ZA8xS0Aj0cP4+Zh
VCtgHXHI11QJQxQNZRTmab4ISWZ8zrG6jO4V0Cwr93WOkRrRBU47xQPEAQJpdc1o
+dCeuZih97Sqznhdp1JcFGO9VqkPSoRT80+gGSk5jdZrssHdHwrIzlA2ex8aFz8m
F0q5yWtAEy59c0isv/gNAigRqHyaWDabZtA+45CnoXoWCPM7n3qRQgMi+sLAsXre
m99Bl06RExz1OO1itVzlfLJ2YiFpwglIAbR/vn44THZcqREZlE73pDLP/Rm11w4D
yWT0kJ5RudJx8YXV9ONrD+UUHrnuwsL0sN4kNdRNB/awTctBFEKQg9ptsd5kPGZD
nH1Bs6prAYzyBjWJEIiMQFc+HgS2tYRSBWcpEtSyxGQWP9t+SuGt7F4MmnSLle13
dOq52U/6tpTzy5yul7hvQLtm0V8L3J8XfEkvAPq65JwGbQh1BPe6sqh6+mM/8GCf
C1k/RizdHMG0o1fhjjIDvtYtERH0FqHCd2kxX483uyve+6L/aRYLAxq2PKiePk7v
/TiKyDjIf4JhpijKYaMB6VYT53ZI+/2oxmppjsAG+cNnJ3LIXiv6yNdClTjvthy8
KyAf5q6nfs3QOJbEmlZ2wEpnkXw7yP4+Ef7CjPi3dYwgHhXROpBKOZ4yRPsl5snA
gSOBfc+AuBaRR3O/4bcoTMUQ4oWW/EMzQv/76g9t3mUgnOHCYhD7Hxa4/zPaNVj2
DguDuzMhCdnafiy/e2ZoHuO/eXDSH2knk80zuU3D6IYsY+X4FhQEOBsvSiDFWR8J
IoBdi+lP/UMeQUX/vxmZRIhRJfT1sT+JwK6P1DkWrO4xI517RS3xs/U63MxtEd/r
BIwqzgFLblgxJwk1V9gByZ3OI9gn5NYuzCy422nmcEWmsGS4lBS7xt+oJYvxa2NA
5BONPNNF306C+37foabcZqw3OIXcrdRR7/q32312fS6D+aXmDsFAsHpomAFPq66q
foY/cFSbmSvGB33t/yA61B9Iz5BvoDUq623NR3yzpLfIfDOR/v0vRJF4Fnsmt8fK
pKtZWXjMVBRoNYUg/ZbAPf1XRcg8ouFdi1TPztJxc/0vkRb0wZNjyFebWiXB6k8W
mEiv5vP7JUljJv8CoMXx1vMHSK32sIC3CnlS2UiQpmoKLLNaXfQgD3smzurktxtH
Q4o0jq7IWK9M+pKXpSDZiU9WwTg7HHndgpVFO73+F98gYs1S5sJ7fdxhFc3ItOw1
xyQ5/gVqege823b3hiPes7cf50NLLQfJ2fFdzrfCHLmnc2j4/aPjk+cLrziIBZzn
2/y8q7JGCHM+GOrl+4d9PcGX8Kb9AWSPL8uVCZVE/AskLzjcVSO2b2AZouic/fjC
sFeS58bLyeEE8SAbpKRt1Z25RbhxqpRLqgV/hUya/0zShZaetVMW4LxybQHclGU5
e/1A81IDwwhAs2j+th8yZB4MyQhjork/XDLz+CQ5wzmNfFNWpJcJ1S6dHCSDkGXB
3WhYBVTzzckcswcTDHPb+/npyS6I+ulXugAElA9o0grJwd02lK/QykMFslT9hs5A
7nIxC+3hYbugJliCQ6Wk7S+8jfUW1f10v8oHdP1F8Q8o1d+JzUUCDcrvTiXCOSlK
bwRNjw5c6LpOO0v+t3ZdqIKaPNRX+mEi2sWXtYwCwBGC+kiNrsSCDH4/C7nWLWMt
R+2yxsH8LvkjgmxYetaN3hbFK0uTpYOb46Wh0bkPEGN+bJkZVDDSGl6AJcMAARWw
4nMF3/uBHuj6xviL1UeGpMH3+0TKAMFXoVxRYNt0uEE0EQ4s8qCyitQ29m4BOCNQ
yF8h0pqI00J9ksxf1sxR4o9/v/5wz3k1aWQFUE1RXLH63p2qUi7CYajDpgGqBglB
NlFSS2zlEbLB36mUZbu1qeF89u6PuBQXdURoTdIJoqn6eGNHC4ZTrlNdubm6sA8d
0fHFHzgbdxaDFj8pBjZKLMDIpvotL8O9D6dLIhsYGASrUepRO4u1G7InWMfK1vKb
YOV0vFTXcGfpzjIES58IDjADKg2rDZJKCI/grfcrvO/CrJfTj6DV4uuCmv3f5SJF
qxBv58rfkSAjwkReSOb6hs7Cwl+YvKGEbmPp/hVSwqocm5DXmf57NQUWFUfUdcIu
iO/xeYsHZ4yli4Hm0YFzz/Bm5OL/Y8hbg7hH6osWy/9BEt9COUMpkeQ/xCiWN1Ni
XDB8iIvw3mv6l4mfx6kVr0/E+MsubFyU660rLVHv9eOz//05HFIEHycTs4fk/PdB
g/vkU1yMnS+UtnxVp0xZ6ItJpYD+xP+WAk+Bo0r1KLtDT0FHdYtFjRkGSH/dITYf
vWB9/W9spSu7t3Yw6u0Dt81rlp2+ZR/BPR3i/ZpeLnKMk2lTfLeBxjtvfcZRqKfz
fjToLwXmeVpnZ39Z84bjF0sB1ajPIdo6xDNslx+AKSfmSFppmm0UBkd9B+YG0Lkz
5cUdNQjqiGgAGCOihy7Mf/XBw1LTdPE/Zg9l01doIVVPlwLzlqmm5hmeZX2MFPj/
sTuox7UkwFMfB3/9YbnX54vwcff2BjiE76/d1b1EqcCTjcqriOpUm1ULzjrKZRfV
hbjwNpNmwO/XezOqcNmFH1gLDyMdVhOFcdfr1FCjfbmUh4ikaQ/I/SZ9C0Sy0q90
O/kF2f16h8JPy2iPTpW4z8xzUhP2MMqpuzGLreMAYZiCWJu1UsXfK43EE/JTHWjC
I05d4TSGF3M0CFQXZIfQipPN8DAntwZvg5FCugTkXV9zr8AWkXnsM313mCm/NM2r
tqrzSR9SpJUqKSmTXwvbUpuPsWp6aTwms5NDHtq/RqSB7sHaIJN/qgvI1hAJa334
jv0lmFo7+AksoCzf2RB7SZP7+Sz0Gn258/wqk3KHv3zB1JSqpFZWtIgRCT9CWD/I
azooT76mgrB7XJLdXTrX3BTQzyRnJAfULmaXgrieQ/uxLiJAYmpca72COXxOTAfJ
/SNX6NFxZZsQwTPPDXL23B6MIRavRtnOrNYzqx/Rq4wiLVRO/wwpTFjmFaXQB0Fv
OzFvx/zFJhinkWa40mnChelQiOzGe2ybJoNscpI5wV1G2FTZtaRb2TEjVx8fVSQ2
WfhwwJB8xLBNNYwxRctulr9VSInjVCiKP3cEMWrbWyBI+P7KuaNJEAN+DefmHWmT
fvdDE8cUpsz0iU7MhXSea7vOjungA6sUzlh52FJMX4ViXXTisnuO05Ua15kIWznT
NPG3aRElw2VwkexTSyWgdbUUHOQ6SnbJCsQvkQLwOCnaFlhgbtGBZ8g4fWD6OonI
NmgcUjDHUqizLA3/8Qc6DEO71O4JE68m50uL2IcbUms09mqkLyxx1qj5r9T3q56L
Q86c93ScO9zMY2EGFvKVox+OLW0XIeIMt1sInnxcfw1nU2J95Wh7k/WvleFXO3wn
bOAHx3Qe56NoxXU4kLEKTbIsn+W34NcUK1+IG32MXMhRqA4Pw3lQF2LauJ6gGlzT
N3z1Xld9KbIGF77l4a1P8buhGlBIMmamvbBqWe4M7vBVfxrtOUEv6beqdtmY1Gye
f51LZDYcyD2drTmCFTeShUpxss1PinYLqa1bREbZL8zkYzB9Lk9ERD+F7B83cWDP
hqxbqoYeQuzJR/AAP2vQYJ5FKednWgxQLFqY91A7sDZvpd0qd9SOiL1wvzR9ELFK
d2fAwLvD4g9Q0XWkodzGZ9oFYDUDrAgFsLnSgITRUHqcft4Ce8f/0py8KeQTt1hI
e8+6kTl08YhTYiPYKpNh3leSGkwE8/zoSNHZh7fqUe6Jl9u5wiRXzNANzb0hsI97
qzk2jFQQL3OaYSjAPn0ZyIOKB8O8z/Q1OL3hM5OHwAuVpiskZqmCHY7dcbengPZk
nJXnTrghHrFxMUK+apJIhwF9CD8BK3Dfe3FBUxHu4XDAC0BGkzVmlpmgLkK4joAf
d6psNDBfvF2iu98FIGF0+qXAf5e1X85gMBn8EQun+jGrkEedh4+hi5f00rth4iWq
9jzb+J8Yf80pBwCVkf/flAi0wXsW5sNW8m/qJMdPSjSeBMIqE2byx+8wi2EUq3mM
DrhMmQZdG/X/tnr6u2kcJ/ECdG2SEaNVH2/F1xCmViGrQsOg7DbfYn2kqGz7tNf9
S/oayYqJpdtFQm74TbB62nHfEgJBZYXq6nKMZ4bSqaMixmMso+kMCJc00t+jSIAT
0TZKyMSfI234MZNSl0j8flqugKVLg9Q/hvOTsExuHWUmRT5WPVLA6VWNcAatipVA
p6SnSEWd72YnaB3l9yCnunHBD9SYXJmJxP+PNweRMLCqiiH2WnSl15vOlVR7NScX
y9c61ar2ZpmfXH7bufuVB39Lg7PzwzZLR9AZLDTtqrMHWlSR4TPxCSGiY0zWOyFu
/2IrZOSJWagMAX/3ZM6ffYe4/ekcfbN1F3ltah0yHuOelu0UtJ0C4s1gUI0zq/c7
sX0tq3cKixrMoVcZ/Opp2zgxFOdOMKB8PnnMV7Mh4cvpBQuJ3Kmk0pxLw/nOIYed
E72fKyuG5Ii8svrO3SYjIe7X2Aysap2vNw/xoWdJ39EWLOyZJWEwwDLVND/defsl
pJs0lv2ByAgEcPGqkNJsB+g9daR2BVHESrQwnkhu469psseXditjh9cwSuWpYxab
+wggf1Lcj6zo9321RkkPsQqjfv5/mjAOESY40p/rCY7Wqhaou3WGOP/H8shUCf2U
Px5sQBkFgNr0DvJg0aoQ5WuFOqyT/43I6QIxkh/FHQBPfJrjYDfO4r5DA5u6HhTu
Zb/VCuv6umnIVmww292s9KmpJJjMoHmt5upb5SL5FmxgSZkO2y8aM8xlbitucDep
IMebbWLPN/R16FEw/UXHkUWlm5z9ncvILxzp+URvAWzwu+Bmtp+CvsCzdpI/cOXL
DzwruqnjnDpwk3fYl3Gt+os4yNQ3PXAqZnf2kMvekUx/pccWfLeP2HJbdUd92l0H
47dvwbRUpS2Zu+X/oa/7ONUq5cn3ffWR2cXJbsIDmD4VU5kbW3+DLKMOZwmUPwxW
v0OYrx8zGrIfw7PywxWvVLn31V3KW3xRfrDGEODEIXtCMan+msQT+Hx6NL9CTrTK
6Sf6YLiCfwT+rJZPIvoAnkwsRNdR3zyysDt7BcbxEytNmPq4Acy5bHL4RgaPn0cu
NbB7mSZmBYDXWk+fWcmxz2muDLsLEd8wqiv7DGWVkrCugS9wO3lqmB1N4gdAtrlV
83TIKBnrNZlGN2l4fCxJxJrBV+xacSMYvZXcaZBE1tPzp6gc9O8CJQn6BLYMdZqY
bugX7hTD/X7Zd+z7/4M6CEpeexV6a7Iv2c+ywGV/5AdDPTXDWlbwngUqEgwOuH7n
1DVIHqcNg35SNLMS1/G7rUBGFcCw5uNqi+oC/snUNi0JTjzwoYIhDzlumNOZdUnv
e8qMuT7UyEnvDPWTfylZDei18mBjXESf7MOoq3/ApVbHmHVSrzk6IlS7W75wadOU
32O/z8k5BaNA+vbO0TFVsF7rSfF3jaMLlWBwDYBenR/Z87qqkqS1ATDLKyVBzk36
do7wemkotAJqRzZQx00I51pK4zMWjq7Y6zyBFxCChiYltIImCxqrKp//zanx9Msr
pZp2V9mSIDwyrmzXkYbvy4QdJaMdamM5eJtkcLgjAQXuPxB1tpBnlO6h3GK8j/8V
fdAVVxC6/HqvXSmO+M/MCI7YgR6kBbwr6U7+JdOHsdcId0TuWl9rTsQcb825JM6V
t/E7NkQ3AKQAFwA1HWV0ezcxbO9HcFTo2GjGwqRI744tbe8br1aGv+EUMFSD893K
dTU9V03FaiGuLJsNzmXjZv2mQahoAf//FS6nZgH4J1VyM9/+tKE5umjSXU6r/A/K
+TXAD+Q8jNdt2UIuG/71x4XxvXM2D6KPTZrMyYEIur0WotWmi0ew4d0Fl3p4pg6K
JgyWN8Dvcww0VF4X/u5bdCMcbwsE8zVLv31i3rDOrvhojLjfn6kuOztgqM9f/4g7
MQd8glOL0RfHok/328yhi0l1b/VDPZpBxNiI2Qz1PxW1QoXTEmCJkrpnyO88Xu2g
PW80bomBUmddjYpqLCGszSTG9C9Rxg7MejQ+n4J4gKCp0NFwpW3p7RE0y1evwVCw
qwhE1B6Rt1Iu0xDB/PU5Km1nmITY2B2gMFQ+QsxgT1xknHtQ4IQGfk/Dgw5DUIiX
Z/eskdnS7nZ6I6rK9nZfMUtwcdkpjzCktzq4ZSsnwmCVHxdbyerTqWc5wtM4jIZZ
CVYP57FjxwcTgDZ0gevQg1/BJAviO5vZMH07UyYqsOA8HgKmF7G7bBjpjOIG9K9F
Z8/aTesJAUW8s7PoYvxKiWBYfL8VivAZWDMLDs15hRAeQlevRNDGf49ZDlbLWek2
ECpdBGJ3h1RMOQOpl/eYbL/a59GIRMWmQQzyDOQfcIBmOTLIoyymOv0LbEiqUSXX
XW8PueI7FO1hF0BjX9iNEphcnr3wWxJkRplQJVNcPCSlXXVHLOhDMoZ7rzD2uZsf
HHQq/OQugTj0mUFmswqA8LvIPkR5/2se7ZN22VwITFhCr80o4AdNh6BQC5eNp+DI
0wrF2+bq6mZjuK08C9uz5Iic0MpnC27h+DlNdsCIoS0zItVu+nSErvGeH/EyXtTM
vyWaTvfBiuQ5ll1ExxeKpv2kKl7RYPSTz8Kba03u1ExCLp/3Za4VNN3KmUMwd1BP
actDt+8TFwjEpeMt6S+JXE3YE9Atp4hMRlkxvjbyUBhyFuTm5pgwwe3KvziaryiI
IO2ABbC+AGKTAN7vjy6fVqwx8kxheLMIl08LmJU7T9M9auqB2g1S5l7w2Nfv/hqm
sluLTEClLpmu31X6wkyXFo7+iBPx8wgbuGFJUOYtLD0JbmOqHGSQmwrplfqx1YwA
VEJIV2OPALaHEWWR8Q4yPSwHYHxQ/hBxIt75m6aAzCyaha/JxP3dNteBZgKe2J1l
2FCdWvdoOSwlxRAc8YAsYkkWDzIxJ89pd17s4IUVu0ynDpTt49RO3XaOZxvXOUO7
gWHx+Ks7g1ZjUcRZyNJW+Xfxg6gYuq5Z1wzAGu5RbHHHlvXHyyYK6zxnsXhC/O3N
ZiZn0jSqdkIdA49sEXa7GjDkHMySliBq70hj2hbUUeEeqgOXKbPFrBvg5azDnyUQ
RyVnf80FkaIJBh8EgURP6q4gv7MlXgJ/Kq0dbWQG8RrN3zILWBHwYGxfv+dX7tSY
6BtJsFgUMNEWdL98+s/eH1hYu9/E3/p8gmOItPlRnboViu03gWerlBvb9FxWsr4q
w/UW6XiGMr5txkhiYNkaH+EJIxpaQfdp01B+/EUINgp2WbYlx4+4hViHKWh0pbWo
LdVUSW3I51CY9XPzBBF/TETWWswjO732sQQRxtyJ0t5rEAsqrpULhtW0N1izI0Uq
+ryEYHdc9GyjbaAT4Xj0BLR0559nrc/HTdlYH1JWFYApt2Cn5Eu2dqeuTRtGq97p
EVFCU+jlqQsZUorSGslvLaQBlh18I1B6vsaPBSXBwSIRxuNskX48oY6JF2ewKQTB
uOrMZKwLgOFQKZQ3LfjlL6YN7E43o9IFoTNb/3ILucwrMc7oA9qaEO3GFECjvRzY
N4O3oVoYSIYgaWjuWM80NyMRQ3/tyvG421WM9hZRqM+VivcwfGKe/Nh38EKM+v+I
WjbFCoiBtr43ATRcn8h01kOz8icaZtt5YzIjVxsG+SnREq5+MGMz38gfzC+eDLod
dhv2ECguG9LY57M6Fdz5DHSt7gfB+OkyRNqGPubww/+v6Km1V3pVk5PgN00f/1Y3
cI2rSyJT9sYxsvo2aGsspSZJLYbR1z+a5Y+HgQKf7ug0hti/azommJAM51TmsX26
UJj3vl0g58O/fgIB+TiJU9RX2LemuGKnOVJoFGQoipbMjZzI7+g4NGms4Px09dqE
zoF929oT1XWLYNrx5fLxvXa41zmCp++Ea4QhLuF6PoyfQu2+j45GBQ3g7MZfLQbM
mKDJ2WuvqKSMT9bHEeesxIN/2KDTNkndEI9VBEB3yImL+mY0dYWPe3dYq/ZZQfAW
7VSpeipi2JMZXWwKKj2WTeEcjqDtIJHpKroFt5mJEo8+LPss/5m0ARiitPVduoUG
wUNnAtUZZFIhBK9ubIC+CZ8kAMrTqhKeBZ6VSa7mKqy9Abus7eYUqmp/KKXPusrq
pnH2xIe8KKLWk1x7DDSlbt8uxcvNKSUN5vDEWxgQBoiqfbRwX2hci5fyTiOYISw8
CBbC/MtKpQJX3yy589iJJOV7mcDI5j/1/oORNXwJwgB9KZGW5tcl6hir7rXdjAlN
JOVuNRcuB7udSJzxzmxNm5ilsOSKN0AA9QjMD0HiyIVvd4PtwoQn9tB//Gswmy/b
vle5/OjPfyPFEX0R1PxO3g+J09XDhs8QMB3QDxs3WEi7pATsW70/9/vdAi4cZdb7
xqkVvBFNad+EcjQ94ebEuP+bpOhwBTH7CaThfhhtjpvknUotdj1/YUYbjBeqKTqF
DAavugWFUla4TaTckYKyMbRqBG+mjUg13ItXzn5LR7hKWbF3ZXevjTScW3MxYAi7
ndh4152zqKRZEcK205K9eIEORpouEjj2ne/SB3yFKMcBRRVpNinJXhL9s80uDvi2
4Xqojtzvv74tqmG+OTLsHO5SOK5D6eVUupIJtBWILPTBWcYNhAEYeGalG+JCwE7P
wxnihMBpHvoQZNBoZbeb4/90gqJDLqha0jV/zXmBQ0IoxFZV0O+XE+ja3NT9eoam
Xnq4skODc5sc4lyLwtxXo1vf8ElXDs16wOCj2ZYrMBZwG9R9prb7f88tq0BHccDz
O3YyinCsZzrbz6Q/nOoYhGFQGzcaH6c7aOFyl7K+a6Sb6sTl5wjmuTvAu1JeWho9
9VEctI3BItT6YWrD5f/8ohsOqhLv1QFWZi5TsNAMcwbO1xDIPLHvxENQd1Bka7MQ
APH2LWvc7lAYmmtJyjjWQDtuix17D3mWEc5HvIpqudqdjVYMJ9Cpp5fZzqK58ILO
4PjBIYVz0SFtXE6PEKu/4jcxuDdDzK0iIUlLB+UGZkFwEYIDyPXPVtghfLcnP6N5
Owos72M8lwT4DaKtklS0XTU3e55ysq7sN00usNhCKC4dG2hZVqLI0tt0IPfw28Is
agDf+b/km31DnOG4BJaPenqfj6l4634XWGmETMHI74oBE9iO24cGqzJQpURnJMbo
NJvUHvGE2siSBx7yZ9FcJ/zUPPBoIdvcXkxsBWs0h7xgjzKlLPxxYj6nOunuopNn
MoUBrxShzeXGa2EhaU8T8BQA80SN4NCm7NKqxTWBEYZJYXn/b8+Wr3Aax5MT1HB5
JwXzckcAWMMaGt+9oUHnKBprovUbT6ZA/P34kwlgGDwZrpY+omnR6OGHcs60JWYJ
0RvbxnI7u4jZmYF6Eax7F0q7oxBwcpxufqWdr7WYLAOvpg1vKchsgEFrER7zxycb
0phVQZC6ud076GB97QQL8Ymtgk7uIpHCdlgz28T5nS6iPDgapQWdkAOZZv0zVWPa
Okg0CcBoS6KnfEh/wldKlSiW45CJiE9w6TpSAWgZeQTM5wXOFH+b2KGIsCvwIPGQ
DUcy0uKuA0RHPoN6w9Ps28My+A55DlQNQUO4LsQmjdkvsdoSSIemEmyxOImP2npL
7271S6IJNc2QS42PMlj8A+9n4hda3VEpldHcLxP0a6/I9ptRgnAybdAXgJWagibk
jBEriwXNu9+vPryA+pETo5LDFYpx3Fd9FzBiKXqTHB/dqGsB2Dk7ucbk2XmDGI0F
irqXGeZ40K18842OCmb2yMYOv+1m33ayQO6Q4tJdm+GXc8We4RniIu4cJvZT5jfK
nZqNsKp5WhpEjVW/s94LldsEytAcXcs6Kp/MtPkLAM+kE1g/SSUs3cjOsWOQd2hV
GzAEINSHOf+CsRKc49PsWJL01wCWi/airaLfC/F2vGZ/bTLhBOLhJATZcsbIXXPJ
GgvD9bhNtKkWWmsvwjxOj0L+zeM6O7aHYw4/fgh8Hw4wFuPheHw+2Otaw+QDVXYh
rsYq3ggQWRb6uL15Sd3tuYl47V0MnFMkpJwdfXlt6XCzijKpnNGEM5UeWtjFqKUJ
y8hh/u5I5URveT2fE0rpN0Y35d4vYmQnFYshztARHPtKe0sWYi4XUg/lDOGAwbXL
mkDXc0SBT2mi0B3g1lKK1JuKHXaKcY6z7nk6xFb/bM7RaFZHOaZJAZudIAXPWCa4
7K6+ZNssiTtlymAKicd7rIIPXKb0w89Yi41c5qHLwAiz54QRRHadYbzhckRaCWug
djXKFRxIhRMOXq69dA3nBw/Rpc03Zcm941ZBldqa2hGwLi0ebRLn4okqD48XJtMA
uB38uoCaHInELgYZ8aHSIN7Bz0gDKteoRc2Zw+juBwKBJlnSs8DEkNeK1+qGxWVk
jIjZGSx6L1mn9uBKvnBSGs8/4f3abOFRybMAZn/aOUYFr0yh9Ci+AmOhf2veaL8j
gMkocHQM1e/RVIGBcmOfkntqFq5NWb4+BG+zBqzpjeCwQ83lzmWy+AtwtmIle1PN
TLRhft1dQxtp9IpraUE7kKX88xzbrAkdGCmDOeBFqrGTn4brt3Snuqv4SIRJRyCs
yGzwu1T/m5ua2XYZ6lgvMNGmzmUwIMKpDhS1bYxo5y2jsHO3yHqMacuIZIxTRk/s
whH9MMXqwh+L5CvI5/iGiTHESlAwEJLR8ZikM8Bcv9RNzrG0edeeJxwlPQ6fqm+2
Vq31aVHcEJ1ibQ8J7QDwZ5bujjgKbv+96oIU/6meaH5Vg+mG672r5pc+VHquAT/t
98rkWH0io5TpKEtZAPp50JjGOaSkj3JBYFKaDSj20Q+A/qY479nPV2hBZqqb6nA9
j0liyXi2aFkdn/i76096s7/x3vQq6DY6Klh8Bb8QL2uLpraDJeEVly02tULvyIbL
ua1jXfcRjPXWCIfy5ZiZXzOKBAxdI2aF0DhyV4+rghaPNz1GGiQE9mCedRAmkzs1
sJkq2e1WeGdKso7adMjO19jREH4BXPAH9bIxw8HL2Jvd9RCWYNKZjtqQuJE0oLko
alOqC1cLC6a/L3Dsn2HAzei77U+sEmSjZulzENyIriqDjMoQriE722CNvWOy4UAo
acvMc1WFmZoyqOxHg7Dc3ymWoiGEaUixwhtKH352dCAws0YvrXUPBKGPn49Kz2jr
0SdM1JTtsPkSQ2hAqv/5xs7KiwOq8BYcXAV8hIN4G9q50Bgu1cMdZG1hzsMjDQn1
nAuHA6VbVCqTSnEol8oBVazL5NpyFlXBkiXgoThpK7oguMfhh6i+tLb9H3wRgS6+
Tii5bmnuyqqdR6FQqnwDsy6jVOWWPLEIBHy8/Y+6CSyVeVJINlfRXw4HJlBZ9AAH
O/1gbKCEGWgHraarzos+4QqMrAiahP4AFz/P9LpoQo5YzL7U93beQuy+o9zkeE1R
4d0SLK3Ykx8VGkQkoISfOWhImre3Asxza7iOL8XK6rQ4jDsSNNeTznXsRi6dzbz/
CyZqrXObjaKnPzQFC2KdHnitd/c16n4K2F4+P+zkpP4Utvg5XKqWgMXR+ZpCfzUS
8qk56tBhtThLX0nPmJi9FGbTBkAZ8DJmX9SLHi9MbggjlhjogKCxRTSjSelckXis
tIaL2vvEXnELgvm3CQFSP3XCf1kVHNsPvyJXQyav4/vz7KgV2rq2YufBIGoh6xMf
gVpYSEvE0ZgoTOlLvcigaeyVphD8ijHi5HkHK3xuWNTFQweMsf7dIjlG1QncJ2eR
g4k8qJhyZULZCaqfKi7Ss14tLoqGTyBZz0cNtjtjiVQf3wPpHp3qLi2fHolO1HY+
kYWZybJy3J7o3nE3F7qKZ4SLg6tyYv+AThlDdNNT/bs2WVPdMpRtlnXhluDW61a9
oB8AJDbzmYp5OSaM7vWYxsOFx7rn8IDMlAqwPpgpDKSjPQpbtA/Mmj32Q3IyZpUE
s1zoP9Saoaz008BpdX1p+XmuVHSnCr2pbwdg5xBgFozDHHLRD/BhXglWyIUMd3EP
yyPMbCtrUSMA3fQCvr6CnMVlGNERvr/QD5TQKac+oU1OjsCLHd2fsLivTV6antOX
HUcRqFfdw56T0NdV59u/TozbwWQlfjdoB8WZI7Jz14QGJLGxGxIkNvqZesWadXvK
Zd6w6Z5Vv/wBaXvvupKoXMby/vX30aC/YTwGAJCaT64w99hW6Q+tU2gMS5x3j+t9
NU75CrvFgS1CtEGZuaBsdefvvt5lQlZX+Ikyu/b55vlnHXkxr+Et5XyGB8y6GfOA
xBFinh5k0w+gW97x6kAeiVTqAbaXj88mEPCymSllYKY7MKK6emHOIlirnkcNDV1/
Zyh61v5/eoJxshEbTnOPPsDm7B8ol+/vQxYaCw8xy26ILYSJpechSHAMo+f9jINm
h6mVM31Y5jo0Lx7LGQhN3b82bXk0P3lBmITmASNz6QSD55dA3mLhsY1JFNOgV151
fftwuTxpaCvO1HN/46XaHme/HwAGJXaqpusrlZIspUbvJR9YG6rIstKIP2+Cmtdf
0riJaGJIK3euH9gnfc+HYUtGX3NIEFUrcrOc3idSYv9o/qec8KVCV65pwUyEmlVN
lphzT7mV7RJg4fRjWiukqaN3FDwOBY5aYAcd2hUfP1WhfuxRXNqbgZ0M5/Cqf1Y/
v9i5G+6Pi/p/vJc7uKw7ucQRRLNXg5/+5UkJ0yN0o65JjI+zeC5H3Yw8kfHk+FL4
uZ4iG5I7EqK90ZgUlfOPotKHha13C7J6a2xmCJMe1QKaleZdkj3afGWGdWSBvesn
JHzCAdk6qPRzMVGKNX9z2YLk2VAAH8hBJJLB69a5VMl0mq+qUwU8O4WfdCkrsExk
rNHZU0YWyFZYksrBxzKZQfSte9UkxUknRgshDHdASXAujBlyxL+2fMfpIdE1COen
VUiTiIdHr8ArUt325YRv+2rlYg7RA1RLThFq0X/7/NF/98VP3e711wfdJBDqrX6S
8DBc556ouk0Fz+HzJxmH5HP5+SUgKIE9BXGoYAS0vf+n81w5Hp/5h3DbcoHx8nwr
dK+WPq6EuNNnhZZ6DTmrzOtSQkREWqcSCkMjwhaknZoUcIvx1eaHOgI2KUjILfah
BypqAGSsN/PtBJJvQb12VFWxyT2rQf9X020GgN3fSVdWzcWFCtK/xJd22p6MPX+S
CaAsZc5K7QNtSOQUbaiGgODCf9NVnOiJDkPNNphiFKvdOv3XTdgzqJ1v4U26uDFL
gG97Xt7rvd5H4CulpGRtQJxYUG22DPyxmx3DPmMbmvwM/hECT2+a3dZ+v3TqICuW
mbcncJj1QPnqUGjbu6b0jbe+fbvG2ycO5gbY9ke5PWxtL3I9O7sEvD8aESYvIzVH
YQU2OxH4L6v+a8NyEMs5a2ly1ij8s+CjsuR/W1u1L6jdKlrkoBFLdAdA5sXWLH3Y
g/1RAoydKEoNm1K8niP3lAFjc92Ktg7LjymOlV75hBNjKjCstVzjDMYId7BCG8cb
xOWLvMZMDoQF1iE9ydcto9IPLe1nnkjaW0v6AckuWBblVQxdtp2IuXeQgWdQtm6b
3yLDGmZJvz9IOtiH2FYqUqdvpH5cYBHiBP2dP2rYSGWy5CjBxxqJ+Brk/oru3MBF
qhL2tbZb0qtksdIaj7p7b8tgr0blvEYiT/9gWEqM+81zDTdd/G4miCQYdAUcHslV
heSBpdY1XSBw8sPx8E/PLcjGZrcjYJ+dM+CJzqFnQIsnnetj1uBUidcGZKY1iX6F
OPkxPuGw/GefgSv5dSCXcru00xHi6ZDM0kAH2UJmnlGx+UaZDfKCXxXh5VwSSKIx
gGi7ZEsLzmefwwsw5s7cskm9wtocuMYHKzJhZuH64h4/a3WcM20I/W2nxgsx1H0j
3xrjTcEq+++YnIxJT17pcUtoAm0xIYhRFijhV0ufMxQZg5BO+LTEvM3Uv8pqpLn1
b+YvEnTp5j+rHpNlBBr15cqzLerXCuLNnZDNHXtf3oV6LTJvtIgI/nmF00zpjJxt
jDnq2A/21t+lvy/fYhzb/LOTfW/B24P03QtkFm1f15YlThqN9xR4hI80thBh3BE2
+dU1qPCSTWBgIM4hG2z9TD9HQSz2cUH8TDuUUYi4tF/SoWzGDb/GuWGoZTVqybCT
Nm+8TnXsmuh2tUsjE8N71Rm+wWvIipTb6djw6LeAKQzAkz1d31Da/mn7Vb0tTRb8
jkszRcujExLMqcb0KLSa3ubyjweyeqOTdMsNBNT8504di+bszd9A4ntTJAE92DxR
qPyOWXHUqiz5i9AzabHydkFOSJvlaKwGO7KSKnwNaKXXDqJxtoDdr1A1QtDV5oxF
H4kPkwtB6iaRWvkalVgJvdAr3jFXZcUYy3S8kXtoyHgFo3z0RTzi4t8bEqmdrkGn
e4IqDsL3TOeNgBQE12HT2x2QsBXLQ+FmHlNoRejgo6zOLhKYdemuW1ddudA0TmQB
BGwwGg9YohWdoLT3Jn7RkghE3q4Bh2sf8keBoyDAjnK3zqRJcWX2D4onc1fkjll0
hBWP4u5Y6ujlZT3xt16/hsxQRIxR/qJWnbSPrICP9vANMSvkGSEK4HlF5Cp648NM
4zOGr2Jjgc0LrQDk8LYArJcasHe42qhGhVi/X4PJqPcUSdiEk+RsPyqrL9VL8AXp
a3Dp+wE8yrptWruQY2Mo+P3Q4FlgNlpUwjp3BHEszGHuvBg4blFQc+mCT8fD91xq
y3d7GuJorO15ikW6N+YE/uhFjoikFOkVZlVRF6bh3rN0/OCqmZ6CqWBjaFLkCMqB
GmxqohFpAkZqhbcV+DERTmF28My/ByH+zwMmT0wSv2P23Dl6Q0rlhIaFuOuBgHsC
KjUnHB+jwrdCNiPgSDiP/R8ViR0EhVo1qlB/Oyjwpmo60woQVJ7YlVi4Wm9gCQRz
o6jL1/xd0DgAKGNEA1c1gzI5yOghHWQV0aBviTfEMjpXWFSoClbP+a0u4HgAFyfb
9en+z02Vzbz0yl7knz2jWNc8DXd94VM5+CsG+ZzrX1uDQ+7WfBQuTalbfka6SlvG
TsnrwQxCv9S4nsgLgUlNhf/So+iFM5E0N+te95yfd8t27rHBCfoFLTzESCuHcC3R
xNwTnZHjDcoZIrEx7lE/K/Y8cOKGImi8Jy1a6JFfvh+aaeQDQqHOh7iB+24U/4/y
VPRstPcGD+CV0/Wz9fJwjiYyCk23NW7XCasqgLcZrDvTfge+/1giHdtOVzQBw5sd
k8UuAs63wiZUdEKoyu8sp8Obcgmc4IvXR/cv9LpW+/nSooM9qP67xbT+0rlgQPj0
I5scEgZMOWfrrhdO6RbWZmdcT/V7AAtIp2xd8ZXFPpBp+SBsgc0HzqOnhjcimT+Q
ZCcftWdkNnT6leLQDeo1hnSQ0J+vf44ojGGx62wpEv4MgC2yZAvkMMioO3fZyNW3
uhfhyLIGCIsKyBvKlqaF7NBc76O969TGPLbNqnz3k8GNrL6I0xH6WJObSGl4DXzG
0WZHJ1ARqqEx7P+PVmybEGiE0kYMMFwgP4qOxjHP+nIx/r7o7bF6xpABc06WvF3a
86WfWXRhg0DF1hJT6w6b15EVw6Ygwh9xWxp+9gVHTDRZgLRAePkPR3QJ3Rj18D3u
XvPW0Srk7j22v9TDE3jxktrObI8g/TCJz6U1jhJfAMVAjO0eYT0O5NrrxZb6VBY8
cC59JvIGNrjuNFwRq1zu6JipFN6G4dAyUbcgGIrR7oQ8eObAFYFm50h1vCptkuJr
byXmsdbdUjMxET0u5Ub+u3ARAOMkp2cKer/fm+FUKB28qD8vGHA4mApG8EXItWIS
z6yI4mLQfBPtDhpH0khJ/ZYujTfCCb/QR6MJCt7wU1WM+ruV/C2xVSgHsQXaXiHZ
786m+eYke1DNJbRkzVvf7BrWiBC2Cq8UpnwYk/slZD3AL0qCvuRfnqIGeSmD9fxu
yOtesS48avCwsIWoWyE+SnkBepItB8nqSLH5H5A1fL0TV3uHw1+h2FevRE/EajBh
ludUW6eoRtmt20oDKS+n85sZhPQC8sVCdG9gm9PVztkWrzKQIAqM2FdLfi8WQOXq
utVvAe/1JmoYPGqohaBV3h1SSW8gN53Q/twTCiL+QbUhCOo2tYJQrjAexmh6bQ8F
wgpJE3VOMXVzb8NTKPySVy1Q5lXlAz/uQ5wZ141GLLhjsNSruRu5IeWwruzESZ9T
CUl7+uP/7aFTNUFirRryZnEHnYQrUYMRCS4yfeiry1dhLjyB/MTbgTkhi2ZeXrij
k0Ju5trc2BpqEyuz7HgWr/0kbqr2ftszOS3OI5zgUj1PFJzfUX280oSkUx7vEHRA
k4O8COjxd6BFzjf4FkNE+KmfK6UNEnXjjphmJjBAgDFCQ6kB/znTRVYTj5r46TwK
sqO0VciUQYhnZTj76J22r15NHXuVUIZBhXp40r3wTGNYdDCm8g0BZqDt//DUYGah
ue5urM3NJEregSStIBYnf4H6XPRImX7nz8QRDB6c6rFd/i23z14BM0KbQqRVhxBO
QWTRx5+n59OZpaggdu53RYb0qShl7cw03HOfmXw+rlVZ7l0VJZzU+7+BXkzEt+p/
DLFv9LB0+VWIA0RC+v/AhwbbyDwTzwzmZkeFFmQyDwlpAWHfItHn22LP5eb04AlW
bThxHfj48djMGdtxXkVjj2D7zkc+H16JBVq+sBhHOO6OErwFmsqdVXmJFaOkFFu3
PV5vw1fkxVM9nH+Hdgpwh8AcCgPChvgjx4LgZPVT9iJkpvjjI0tkXCzhrVFrvdkl
uWV4UtFwFjlaJW3S2Zj5hM14lbOxaF1GzhUGued1byUofbCCvHyxMG1hNjCYjo8I
3eWWnS4QekMbi8QWq5KrcDe0I2Is6zoNIa6TLJ4aVufHuTR9WtvzyMTT+lifUBmr
IcDx8zpTbdgxl3AIbG41ZT062v+t2tXQ2XgFLhDVX9md41sWmylmd0WZLDEFNkeP
ohgj1eCARC4GlYysgFC6VcGkBfgVBmFOTKsaJWrOFbMJNnWhScqkOOgrbpFQIEi8
DY89Aw3TYwH5qrxh927XCnYspO64furBSIdbrTgLPlSjb5yTqIWbjqVDLa90bo95
74JTtb2DTIBlcVVEvGZhPI5ATvRg7vv+oGaeBeIlrLDU+qJoNbWn3z+7PZxFrAN7
63oewkeRcuuwFgX8hi8uZXkggWUeTx9TRK252P6IKezlPlK2FRlmGaCoOuAQf+et
4T6f4gZJobb5slg3+P9IvQ+4HYteRmRqDklWXxAT8Wi/KBsdNDSOUg3rIU+MBUdh
dF8inInolfXz8mzS0elq6gPcQWbZct9e8HVpY7/2kligHhU7zlYyD5VOha0NmOPH
8woAnOKkL6oLmmE7ZUlPJh7YbChxkfz8WbsnGFt4DvQ/Qe9bbZW+kz6OkHD2b652
62qBSMlQiHEOmwptBZ6DUsgus3iC1+LQFG6oQl0yNOjF7nYiUDuMztxIgW+loVfZ
ThNrk0oJgbCjL7QqzuHwXRdqB2ddosSQRqpANs7qBX8JS+kUF+kLiuI6Ude7A34b
xFQ0zmnrPh22YSsOueMPg1KsLgGgALMT9KMDIh7kxo6Il5E9q/xU3gjIZumc2VxQ
Pf+D1dDdisSPYld5vMf8Z/iUDzZZVgYMd0VSRU3/t+aqHcp6jf4Ec15v7K4Q1Pms
6/YgdVc037cMOOAJ7KHDt0Ib79XMZs010Wr/TnnBHVJWsRow+mggNsGaoNyqD8xe
Y7Ohu1kWwEjXcpTPvV9xQtMddTSFe1wm8VwjMwVifQMsMFpfpmao0qqplEZngs3H
Ibr8lUEIQQkEJjKzHydByvD4QECeuzP3Aiso21BEBuDCd8DBcWHRqWkvc591S11p
sC02ZDJofBvgAp+SmAy6l52ZSBGNuevbYr/7ofo97SSc/orWG2Rc8Q3dFoLYYED+
M7MgkrhRkmeeHMSBAR6xM5G6ioFBuHADM4dCVK65NXKTyINhOh8bDJnx7x51Xo4/
K6yJXb5RL4y42h0U75movi9p6TQVZzlZBJwzTSMuXLFJIN1PSgeT2hWFLgauW9Ja
rKREDyi7rkpb1Bu2gAtRGfuNvetglrxx3CLvOO3HnSiMQC8ygC4POea7E5cqy3J5
gkkoHNHYj+y2m7GUfyEbf9QArm3dXNw4iSxtZ33KPsakqbJhvzErivziuNIdcaxc
u38+OjciK6dwWBhcGB0Mstbn9nx6EYriickXG0GT1kgxpeMZg16SXnD1NROSgwzW
C46jmGLBnmQOZWihvdqoPG5uCanLaUcq5LI/1nlyVDfFFqJ0v5lc8oRxDA3kasjL
K+BmOYPKa+79YzfpJbCzbXU7btAlvSLtWrIt/kviUWit/wdpj3HQdHwjmDpAc29D
aEFZAi7d3pvnM8bX58/IFLNY69L8daZ0ITKaSUJnShJSTa6usv3vNMb/t5i49oQd
IUpeOEjower+kP9Al7pPdw3TIPE1IbXxqgQtOwnrf9P+xuevdzBEnkaNzczT22Z5
k31ZW1ialZoMZRZtq1N0R+T5TmSd5RLt9X0QLn3dgADyQsdxq/GmMf6N29YCfTmc
M7Dj6sDkyaP+eIYeuWsonfnGrH2NsrVX5y1gF1gC6lLwWqOYuPIkspzi/8q4LK6X
ebHWx8A5luIn/D9Xy4Te8H1mDZoHhEJxPKxru9BWyCsnRE9EXIQMI6KVOPaIPzYL
ibKbkWOzRvLHU5Y79fw/kfxoRxFD+pdZch1EGm1U1OHIy9eV+Eb5AnqMLJXgbq+R
JjlsbYyQmHXFkLXoCuazKjgExVScShzRMk+XdJuukRk2CXvVSFEk6+KwALsy3bax
UZ4bbyvuKXqskzVnOmlh6xlomKGC6GU7LT6OTJP+bPU/Y8hIHHlHIyIhk9mdguCx
4JdGmBlM9Hp+qA6RbgEFk81JPYFtfuwAGbE2K5igQ0AebAv/cFKsBGqXbZB+84yP
K4Z2sBSu7b8IkzBCdPk0q+ptC844W+2nLE/3FQA4P6lY1ZRIwny2luGinh/M/TGX
Gyk8t6ePRVAHp64Q1ELcUQ32WOgd/oidRLtjP86UtCbLKSXEv/Kdt7Ze84Oa4kSw
75G+6BRqANCeQcYh1h8rfYoJnvkkqP/bqM3Jfxr/Vhs2eMyfTjHd2/YHyG450EZX
vn1E6BzY24Ot7C9MGwE/x4wn6lEAXWC3V0g5oKVLBYz3Tnw3/U66MTtHMvwjMbDn
5LmTznNw2K5tCBom7QdejJ1SIQyAvTAkSoYDIhdT7bGjrGo2/pOdhTsMPaLYY0ZJ
KWgyRXi/TXd/D9w1L1Ok6gBWapUZbdJiqzVsda5cDhPUzwKMIVxgawi9qkez2vLc
GY55w6KxJxHKzSWmXhTS1mVL6eVmVEh+LVHWZbQ+LGy+ojMK3YRFez5vBk2Tx0Nm
buTgpSwMhswze/IyPfhiq2FZEV9Z63zlJ4kBSrVMWX8XPPve5tIcvolSeaGS5gEh
5+UhXV0Nn97FiZ7XmJf2I5152ECc5f5Wdq8ErMEvUy1PnAMySFM9TC7Zv2EvN7Hb
pF/HLgFm8q9sMeCrjbBj7Ed5H6h0gPet00CGvT5s4/X8UyhR9a7pQm2fHvs9CwSJ
7trt8y5J92hLOslntjqJEhkgJpHIcEDPbezyiMXaihdDjfMn13f7YFFqK6b7x7M6
Hi8fPgHd3U/jNTi5euDuacNgKyZ+1T58m6zwC8NffaW/Q4CesoRyamYbxQRtbweH
gBLJUNEhrJlk7259hHk2ZhXuRXL6gBel0juNqeJ9QTIs0sum5sDbehfuNWzxyuKR
wU079ZlTgPCz18HGrS52OqCd6zPvMwa/q/Lcfe0WJORraBB6YPUa+tQvQaB1akML
+v1F7XPViwNC5xvxmMRTOEKjBtBISY46Xz4e+iRlizW4X5eeLP/6eMSn3GJ5Glor
zzKxGKPMZTXnXKETW4XVMieVbiorEfTsATtM516iVCDPBYLSIWqcU2uNMKYFP7HY
kV7Y85LTnntSn/oAC6ocz9d7CSZP+k9+f2Z0Rn7NVnwjodKDIF/eHbJ6/kC5HQik
GipsRfK7RBXPAZ5iInBuc9gllR6xcDG2w91QFF0cayW4R/9AjuYHMNCjLrwl3idX
Te91VzorwJn1FlrzjBxfVTWapI+mf1ytnEyNFanf3alH5NGFwVBzepgtlhOjDKpd
X6PYXdvZRVzArVsmGGknY91n7WUPTbuKFJF8NKaNtmvr0JdcydbFlVUu7qXSUn8r
+s4cvo3vrOt4X1uoatPzgoPD4XXHd6qEin0setYqYkJptKEiFUPpN92Yiblq336b
RBiYOxllU+T9dCk/c+OGshHQcGaY2LrJHZYixDlHrYM0bADnRjKUQwvBTmFnWTIz
EBIDUP8iWPTo0Xn6UEnnzeHbaQdYnZg/rkcZdYE0kT484ghUxDfPSlU7WP3wC37N
KTyRM+24poK+CGiaa/ADIfIjJqv07DILkmdxWQlxmd8MiIzcIFXgOkfAto5a3cuA
xcB4rHW09+oIXzY+UJUcm2xAJnN+K06XAKstov3H2X40J1osfL0VUDoS+LET/5J7
l8V36kQBTDTG003uQwKTU/cj28pMZsC2Uj1N7CgLp6I8yRlttLq62X0jZ588R51x
2fCbDVoSs62ge7dTXABESCbWiIv4g6+f68OBkIX+PSKXUP3+xjMiFIEpsqU+07BA
JOIDyJE3MAzHABK4pQHojsWmB6vFqq/x/xvCHcGDS4mqUST5C5QymAZ5zzaTzW/w
Hp6drWo+O3IyuniP0oXE02m15PGQVVlSLiCCbC8rx+74LzhRBRUlUc4hKMxx7KXJ
BVEC1KPTO5uww5BfdPjxm7wbAXsDs6xHLnAwrlZ4ParK49ms9J8i52N6+kaeFahe
48Bj7CJjfD7uGTernc6t6cKNKomKoYbDpdYuNXGlQxHEhqVdII11cRF/aAXzuM3t
PFU+ueJ14GoCPryRScTJ/8PGsq9mTR7kvg2gkiM7y9X9HZDqf4UpBgJFLY9RDfSR
ye+wR25ex/yvMNGRpbSaqnDt4m4qUPpvN5ijK4W8PO4tdBQiRUAfTDkmqdo373Vw
FSARz76YzX+OS16Qd+oG4Nnbr8vymKZ5NDvv3zSMP84mD849s0xa5yf4vAhS9EOl
ql38dn+d1hRkVydCMs88ZU62seQlHq1ePuRsY1hbV2zNSaDATxuGXMPldy+FXqDk
0f7cIUz22jhAN4kQY7zQ61RaMwdHWGgiQeo2gPqPuAlsvQY1k7eq1SHpUMgAhsje
iShOOtcz2qYpK8dTVYsPipwanZu/+nfC2q0C6pflOuIrLbt9kmulcPBfotWnqhfq
GcT/BrcKBw3W4RtE7dW4pNsqtckimoz4rdLvaMI28igsAEjFK3+u+RYQRsa0hP1f
stRKyQmC1a/jQ8+4oE+RgH/nd4A4ybuWhOtOi2SIvA2K4Ttm8iRWYWJWeDZGFF6y
rSixYPH3hkMlYzSLjETqJUVQ9jnB+a3cU66pJmhfz0oLH7NhXRk0KiolS6qq4C3j
H+1q2isj3O210/Q5tIr+CAqRcjzSDIjVAYCw46QEunP7g8bEs3MRm/xqjOlg9Xqq
ASpitghLtlmHLLhB6chCGgYpLNi7+RKyBoHORjdv+nLwsWquGXWPk8iD/NWn81m7
Shw1rvJPnwU/2MFB0XhyYJh7sR9DQK4FiijZ4gbml31Ou527nBbUVtMwf020YfrE
OJMmm+VYlxSZpQDKFAqJN7wRNQi8SZ8ln1Ne7WlM5U7I2TKAB2VbKW9ODMn7YDI9
7VQ9f+9YKpGLcYtBUEXWvp6tI2cV+EQXyCAmKLZjymqM/ChZOGblppcwdZ7nHHTP
4FbcwFJWXPGFQjD9A5e+tbQckGrAO9njAd1+seS7lM15WFzSW5hTmfoehgj1tdBx
M/eovhQZ78hSdVoSJanMxz+niacR01i93XCVr/Rv5gguhwEumDNQDy9IaR3Q6Qbv
WmfJJ8g71pUpAZDEEv2IFz0lQIkPekc2WN5ewppZSh/PkSdlThNXruj73rxOPMiA
ATIKsH1NSa+xrboWg8LPCEBwUTzXx5jbxsZURz+ekHfxYTwvnK3bqDKCYYJheBg/
SXbH1NF9wstW5OxCzsANRi9Mj5PJhuLympMc+WIQDdlLg/avPWoyKkfKLPcarPvh
DeGUO/abW+ajNfDIdJ3kvwUEnggjfzK5nT/iPWSlPMXwMwdhIHIjW3qEjy3KchCS
khNs9DdenEGkNDvFhVC0702Xym6iI8D15Vo1EI9is6sW9BFAE0OGtlvUTKBml4dt
O/tjviMJvBAzWU3R55I7Jp2G1TuDN417HVq3rfnVP5aUTn5z0NL9qdA1pwf72Q02
GahpfziDQNuoEwmOAmSDKpRSvMqhl0fSYTP8X8tqaOObfg48qEKD0Y4Eu27NEYXs
Y7WABkWZwC5fKXiOgVCn/+3Uriis08YRB+Ssg2OCyRLoXsRmLDqV3gelevHLUe7n
IaeND3fey86Fu0IFPoiK4tcbb+v6r8+eCDS/vCexCu0cp+dAdAmUbyxAoH5PKNET
/Z8vmYWh56C4MGrgAw45IgF9cbVzWCaSMNnmfD1qS2xC/3enAA77fNSCscklcN7/
LzAKzth6n3Q9J1osPpYKozmkzUslx2Ih8hyC+jYszA1ThjkQ7Dwa6EQ6IAP5wa+s
BIh1ilqHug5ftfsoFHX9naEcXI+pLe2wS2UOCaOsKrGiBMwRTzvpToWCNnva9Wn/
sXqHXwyUBtAscAxanWfJvA6KS/i1fdtZ649ci/qnzJ5+C4QlEmBNLNaNJOSRG+Lz
EFTEpnLtfgyu+mOV6hlTYOP6uM1ZuBUdefDsvEhzCLRrARz/wmb7rvXGEojHME/H
tImkVIbekG3ps2Ymne5uhbBzBaHqqs7+ngEPO+ADwi+T0q9nzW492kO9FSfS9zEd
ahzmZbAZXWQwx3cGBvK4LY2zs4V+1aa6kKXHd8EG2KNqoudULBA5HMC8Di7Rmwz5
y9IgIFPQ9hhMQfrs5dEgvcMY1hSOEBm3unW4zuB3Bgr7cdOuYWX9v8+DPUkc1Ghn
1Z3AYNsJJGGTgVOS9UYQQtAGoRYDW8cWFPyKRDMfRQvBtUMlH/L2lDhFyES12P0b
JYBihQg/6RaK7Wf+gHouOrbBrM1SrVjZ99lE5uV95bnLO8+5Vc3gwXTjIJDqn6gz
GgnolhbkAD+hDUP3cal73wxPWjG/EPs1g1NtDGOgE7sc2JeQ+6xp4LnKtcalMY9o
CjG1Sz9qKw9XSfZGh1SYQFGXLcQr5exaKb00S78VMD7FG/3l0tnrprn+tQhhlT0l
rlCNMSgjSACBo4NJFCafMGdwJgXrm9p8RVhJUQzUr0a9nikgFwgz7NqI7x+f4LDt
nEiY2X4gudrJC1+59V9or/8SVuVFqj/yttLiWV5zIleFJo1GY0xp897gsfBXqKLK
cX9nLSvLvZ1gLI/jxFZJofmqMJsvxpYNEdlYPnQPvO2Kx4kegjUUwrlzSNTx56D8
xhLFvMCcQSHqMLLlgC7Od6oPO2vcBzL9JILUqzc4YG6/tW91pYG27cnOE+46XtMB
ypn/ou73urh7/rHd6fqGEwc/MrHmiKh34NFyzt4ODPbEzRlvK9Oi3Fd2eN2EnWnm
UayOR5fkCccEHqrkIQQLCVcwLLee6jGkC+04kVo8h+7ybleEo3O/D4DzzvMI6XJO
KVCBZA1JJVSw7Sh1k/Y7jw6PMAnJWBKkmcbDRhGE7EcgcKruTqQGILA0I4Oy8/is
VVNIN0PgPKY17C1enBVLlOf7REdpbyHAPJDD424sklO9fL7+ABfkXae3+gRyI10Z
vWwkerFLveefkm2Jbeoqyw81sL2IgAI/sJ2nj9UHZ4atR9FVOwxfKOivYqTqRKqf
1SeQnoTtgn6ehBYEWHxsUNOeEFNwVDjamfcpBQaNBP6+8jdey29CGUnW+bE816gn
YcQ9U+z4k1MwfhZlyaWbgLKlLxxvJPePji603SLungJxHEKwf54bL7QpZN77JRwy
jRNLlv6LhzIo+cG0tw3PfRsrSjK6DG0YU5+ko9tOnny0yIggF1SmtOp5j9r12AKD
INcnAmaOXiQFJZx/959aBZn43UTVkKXKTTuBU2wSCjzPpFpeW0EZqZdiicvAA43I
/E0YikKGF1rHYV10AHLgPr4eMOBBcKlPxjTOwXZ3wmoC9i4LYz61NoGt2e54TW9h
qcQ8gR0Rczt8AeU9UYlGdxGhJMAdLMRnyFeHTb7MQRF8HDZ/TGWf7f6IParKpYof
OpURl5XUTihBNlFGvJUuS1DSQD7ugIn2KWjaRW7kB21CqKUtNa9PhVR08HYZj468
0bSSIc4bCJcsoC32x0BKRxYwa1S9Lu3wSVOj7mkCg5vx99vCUCxdLBjJnGmfveUg
uP9ra4cN6DuaxDTN72hXMIez4PeTXRL0Gq+y2YCOSKDphNc9+4yaOQZY0guEOvhw
JfTXaMlUjpReBpT/4pCqGWsYvdG3DSNxeyreWvi85pD0DwLzptbn59mdThHnWWl+
sHphscv+seY1r8U+y0pTVbE1/VHSes2J6fw7k0BhIiR2K2Uqn9DXAzOzBv5H2pTe
0mbAExPtJJE5iwGq8OGwyvwZB//9d4UAK5F8KfKvatDkl3qCdVyf8lLWx01rhJUi
M5QRIZrs7+hDY+ksSv+XNVpM4NgLBsjanl9l/vT8gLfc1jz4qRwj61VWB2kLpU5F
8SkFBrQuGLYfhgl+2fcsFI9LUp9aMZMUOTc5SHmz6M3MygzJ4a6isrfrUSYSapGs
/SWHYj56ld8V/N06Zej+qkR3lR+Maw7wynvJX5p8vbzH2u6xjIh7LjauekFDmJSH
1pQ4zWY/NInm9rFdbLx6j2e/44Q1o4gLUZnVkFbSCcKh36vDZ0mo+B7jwCF1IKDi
leef72eG3B3QHn0op7HzXbavTizYtE89dsd1ePzBCtVONkLbVPvypAtKbGe72snv
YozTnG8AoeLNOGBi53JVyC6ZzM9tjc0G7ZCX0mu5g5szyYRMK5lJd/GSxKZLGYZI
zZHp72koQD42taNefQyrGiQl88b136g6ITulimBB2cqjqL7SHVhEscAcYiJ6cxum
/h5oUETNmGOJf6EEDRq3tSx/vhLtWYpNzOu4pWgKggirVPxcBfyqQvHmshAjQ1+k
6Kr1TqlhJe4OcSNB6cdVAhrVVd52YhiKX6uIfVoh8p48lIjbk9u4hiHWJBmgjz0N
WT7BXVXN40x+sWw9VsqRhVyhJ5eWagOhCA6BJOr7LkNGjLHI682CEjSBVsWXEv+E
7PMPyrK8/RinzK8RlbEKxo7gUxmD/J2o6/9T7t3WU6T0j8+wMR5FPCSpP9r8paYB
QhIcQWyrAhsIEqj3lJMiNLxfvRjM0tVta4nFpKdxo9laBADLe2iaqCh34KlyEhes
/ZFQgnD4L226deQOiejlYIu4fUt/7G4K5/lIRGNh9JE8+nihuxEYFVUKjZvvgFNQ
5bblHVw2aHAlMkq6Hmq3YNOAJMjMoFH305pMZqfeaOQC/bOJIg6LUpqL03Gib5Pk
HGmoArCyOZ6lTBWyghu7j0l4002v+8kKnNxpfzATOPSZ8T001eLvxoSYyP1Z1QJm
9m6G7lN4gdQF9LeDclkPY5P/JgyY9dTzxF2Ub5iPbQCNlBX4Jkx1Uepe0yBPkuy0
7MVcaX1E7/HfL2mf/x09CdgpKzQBeS4H5iT80rQlFAD/yEJylti9y1Z7N4mmdZ/h
RCBZCNdIW/sgz24IJ89YAboZOEEGu+gsphoNLKFpH13Ht1btuxYVisN4Q7jW+HNh
O/baE8pWr3BNCkHNOPKk8DmZ52KiaHI2bT+N5E1gUB72EW9a93Y4JMhtEmePe3UY
JDBqDMGHPifym6azYdaaZnUtMk/RemqjtcUWcHCnhBXn+A54EblM5KowLUDxQT80
vHb/McQmfV/jtZMKz4kht9svRFoJsY3uFFyrp6S/VTArzCFadbqgOUvJsCAfM/Mi
4MgCNuvaGqDNE6PgFBf1rNGNCVOhG+SJPeZlizvFm3LwcGXdOxpNkF6ChFCgHe/5
JJm3RPkQnlkMJakObqScyECkGdBHTHM6hQQfu/7vImNovkdtaU2mQB3k+BRTyY/Q
DLT7OuTNdnLwu0FyzVLXsIjXQCKwSc6ip4AbzQ4lwW13glQ4Ys0Bzq4wY2xAGW2y
SQS+G+0ubpWFk02DPHAn/abzkj0VKdKBlJPta152F41VKGGSnUWrrxu7H9shSAu+
CAvP4W8svfWrSYMHwyqqo5v9GioabeAipIY/PwzXayEJyE6au8cYWBMVsGe3hiP7
0zzp6+fMHYGDkTg70PUuA7iA6imZvJgaR0dd3fZLL+VUig4tYnK0mCry4RX1Ojby
K3JdFdHMuQqNqa0jB0MbLMo4E0rlFXHudaivlakSxqtQJZaroGRGJ8gpn9Bb6bSC
EAikydclqlA+m9JM/4Vh/mCrSs7M558SRaYto+xqO4s5oOGIStlwkNvz/66JL5jA
sp0e6EuWEVdJl4oQJBmtz6Z1K9XPBgHrWwt6vnMd46mHk1UNZoClAQjh8VQI1hrC
eTQcWwxM4OiI3i4QJ48xqoHt1FVmobj1QM1vMNwEI9E8k4jQWE6LYSqCsvMj58LF
6l0kfA72Dk5GPrH55Ad50uJ3YQw8q2CVjjBULJhJcXKhndxbNGA2vEQ2EiiRvWFI
WDVjg5llFFiRUg4jpwU0eF44QraT9ZmZmkfw+AGono40cxqb5dqb9qH8p3+5WyCA
LmQY/NSG2dJcV1nI5qZfS4zVvpabcDzA6wYmwXUqFy8bsqvVRI5RaN5499qWjFGn
jYY3pfC9C6cR1OiP8bqBTVW8JV1VanQibkbCcMz9aMf9X+mvzrVgiTdHndhvUFnM
0OjrBhLYu2Ab0ZV/yivlzvkfJPJg/Zw3wzd9Wj0S0uJjsKn0rgyH3K/dCf40wE5v
KxzwmcSucjNjM0Y81HOzuuFqWuBqkNQBr0b7XBD5cfHQj5NfinKRez3V61u84kf0
dUVApGjfPHQQyH016wh8zlzI0mggOIMSGsJbIdDiCKOkrBZnkdOGQlWyOLAXSLMZ
aeZYqEPcvZoHHX1vxzy8lFkibN6zA5BzMTWX+Y0TPnFE01wDZh4ny/ZC88auEHhP
iYl/j3uYdgP9q40rbZqpm6yje5V2TTjrx29NRCnRAVmvLLanMSEjygNhvTTqan4L
s+0oFFfPTqLGKF7ZB9PuGOSd8WmmCWfyKRkNQMbZCzhWX2GQ3YAp3qqNEG2ze6MV
E7XWCeD5dUfOlQ4NHwX51EdM+P2BF882ov/nhjGeLpwdZSYDSeDwYIRtDuImKxyV
amGUDRZX4abZaVW+b69rudL2OoIq6KIvQKSPGxGXwn4edq0HBh4S+xbXjpqKLobH
3YW7DR/FuDpXTMn1jECYWxol4Ip3F0t/zcegjvxalsU9ol9y+qf/aVoFp+AU8RL9
gFO202edKaOF52Pw95dqW0dxldtLFfEKQjuM/btuK8uqjpYYjq+ztZsgN+l4olMo
hLA1wafBA5LAES41QHWckJoMpRn4tqVCEuM6j6FEkApuV4CXp1L+c9h5Kyouul1k
nbtzm5vZKFnH0rM1lObwNLD/Tk7ILGel6tGtumEnifbangBNNNImCbRzXNvLWPku
niSVEBJoK++5qhRWGtn9UJ/HeaoWoJTSThpMfo/eU7mLKuo6HjcFILvsE3slml03
1cLNCBEsKSyRYWeH2GdV0RuHamqAEXGu1S+98wSil3cL/O4SusjFfsNQ3cVF5pw1
pYNCDW9C1Um08/Hekx8+U9YaXJlLot2NF2tsExgt3XcPGaKbYkK3Mltd4+A3GnLk
ZiFmf2x6u5z9g8QFfOxMz7FJPp1weiscOvJID1oVhjxmZzXsBul9bGpgqM9Nwe8D
OCBHZ6j2rbcGAGkdQViYSazXN6057W2kH70dq1LdWeKpTAWN2QTF0uYeKWupwprj
O0gQAYY+YfgoFEs9l/qUTdatZpNxegjwFClyeCzRgU8LoPOzCJTgUBkLVI52J7PL
oloalV2ONS+RzRo/tk+3t/wGqCA59us01vRN2Z2rMuN9TIXsMQLg/dgCq/TxylOu
BqJsJ9+7j1YMWsCSac3hMqYdWCAGSf1Tpu5BT3yu55bcHRnr72BQMMc3a8R+0cK9
CsrlbVhMzB7tYj3ASovtkS7Aw2ZnnddRlyZCbt4MBIans2a7fgM7ikEWZ+ft53hs
/Oi6E3cDx9vH7NFlttR68M9U55H0svWIqK/Jhyrrt3ciEyTMmVAs9dC3/77KaUoR
G49hqdjK42F7KyZE9Etqn3sbpQuGxpRbUwij34QIa3UhoZzsEohb0LvHegoYV97J
n5cZHNevZ8SLIccIKqDnH+zKUxDMXsDkekY1U+TDwhVX1e4MHDTg+MBp/xhvKvoR
9WtNERKuu3H24yJOM+COKCHZcvowXD/2kBIs3ILdVv1IW107GEL5nRQhhCnR1hwn
0r0ODA9XaqXQRh2ErFKOKtwS8SDEGDNDH2IKxrc5X4XA/VXVdZV323Qw99L8R8Nr
yJwlUZIYRISL8J4jpPxJNJ8RfSxtha/8c5FdEF5zmaWaUcAmEnzxDe73MEML5vff
cWJnOtmkZBoT2hzbjJXde1MKbZmnXqJiBKHeaI7BkQZzAGunQ0Im++3W/6/57OmY
KQZyoN0oL/74aB9oyPI0Fxs0a3ZOZc27A/Z6JQ/3UtUNJ69eXFqqhvHY8rkFMztx
eLkJPgsgYEDF416Cej9NShGh5S2yTREeVwtQwXh9FschlP7Ez+TtVMjKg/nRIqtR
nK79RKkMSXOCrOSmE97iQQXFPX5wY1Is2DR4nlbSO2CHeoCmJgV/fiTm2w6DrMDs
b5bWsA2UYI82Jxb6ksM3eKFSnmcax0Xkb0C8kJtPL/O/hWDyoQ88RBBrjhmWYMRe
8F0Rl4P+rS4e1u/TuNhRQG+Azx1clq32UqkV2HNAXyPqrlkLzL2TWe5shZQyFTBW
IqJ7iYLoEprWM2TQryQVXSDY1mi+5AkcoUSnLJMhw29jc5huqHdlmPA4Qf4QEiTu
u7yzsbh6/g955GEbik8SpTALJyNEaIGq7KhE+x+E1NtOy+iussWqM7gQiHSsuk3o
KSXPN9ZpOwmOy8f6j3IaxQ3K8sYpRS5Hl1+jmAkqc4AUxICLai8ShyHtE/9hdL/2
+/3x5QodzMiyOW9JJ5HdNH/hOgSAjWd2e1Kf99dOUtftYSBWRSExu2m/ZSh3Qumr
war9wYFLs9lWgzjMRJ3eBq6F1h3KcN8fhBmF7fHxbqSJX8fM2aSH5WRlbyL7zWns
biSv58zHEMG1iOcF6NEkbi1tuILcUQpRpO/AWoXPeJmT5GMfNXLHC7zN40e2uJHT
Teemi2Jlk7I/ylOgFg3KzVYXS+Xi+RNhhJ/mpJn2TDhKxdbkXGXZsXRwAl/1qsxg
OZHfiNqrJSOJm6pzHVrrBXBwbUF69th634HfGay0daW0aWHZsO8RNLtMvgCCe88o
c4RzPIJgmWnyEEoIj92lFXGUHOFRqhX15wgQX0kCqsD3ZDLtMhaQjnAMDO8CpkLb
e0uGy6hjLFM4CoZ+ul0v5aDMvrMwUudro1+1VFg6qP29cByKtFITlqM/s8CsSLLR
8kBG/ppDxc/XH04+p9xrflEtbFO4yixH4tdomJtkj1gJ+qQ7h94izr2vqB3BoVv5
F+WjbNuiB6knzFuBkFeLHC1TRE5DMIfzLmeAbRoX5KgRa8EBazjJvtM4GVorZ7FH
kTk2SBwaJC0gEyGlg3apOOyOvj1uPBFdGC+5uy3CMQeOIE994Kqx9WT8bIQspolL
dl0kPzTrORAPHMjR6T703BEvgKT3AWBg4Ao0ZbgVTQYeqQPzawcjHJTZnRkej7uh
RBtW/xS4d9SRY4uSrKuH0CtrnhycSNs4fBRQnaX1ruzWeEhnQPu6PzSBDITSoy5K
uNWUF4P2bbbzv1lv2Fl1Pymy/7RPx4/8a2KPfeGZ6PMmAowauu1jt/uWzDAQ5odb
wz7JEl6MtSc5d2bXRcdlHEEUeZl+9eUu82IsU6ntT9gbJAuHzWT/VAuMenXBsJX0
WOg8fLS2JgIqk3MErbQ4RHAi3eQY86cXagoZwfyNgNikY17oWj98T3/A3zXpR+T4
E4G10XEzyGrnYNCjBU99xdLOP6dhHEECQbFKiynBcaTo8KT6rnnyJnSsAsDNDI0S
k+KGtPmDlc3jwDJ/6RiO4zm8vL1TjwiGKBRakN/zmXsYED8fOO9LANfahmZ0VNDG
Yt42yvNVJb0nlzhq7fj/BPYvjiSXuY2YPCYQ7BZWmrLFvHfxFGl/SZ7/QLRJ5/jX
X7F+HhjgGw9OV4tu+4t3fAJ2rrRNctnS+amnoeaf15SAhf4qhBSLPOW79jC4rMSa
S+pPzmV/jZqU/daaaZlkPuH7/aOA3pda1gzfgWSLYsjFBz82L4kfXMlFpxDHklDu
380PgikeaO8l77FML/dsrQxtwV4bjIaG/4L2JnBAUcCO8RNevZGaZFnYB7Rx9I6u
gmSh45TmmvN/3Ty2x8I7E5yJaGTln4GE34tfSsSAusJqCzk+ttpLmgrWkvU46RTT
MKPsy6iagYnjptquNV2pzWXizNp1CoOyHTrVpuQU14tUubyPoKyGQw531povLBar
SQbGIFOL8if/DXuGwViIDAEBgjhwBsKvCZv72RWACLIvwzuKovWI/UA9hvBaUjtl
7m3i5+k0C88Mw72v3Vktt2TtOfAeEQ0e2EAy5gKkDlckBTVUwhlayxzM6iVv6eRn
9+IxE+paXSvRs0O9liLSbv32Orpjv9fx0N3HvlZxRzCrOnT2hDEqLfkrDYm3Jgro
WkhAZXh7nJt35CHggRvnW25ZdtQv8Z+k9NA+8TZeORBNHDHxaBsXDptGaBhL0qSw
eO+9S1LFp46lGvVYFTZeu/fqUFsjdnhe/Wr8dI88jax2dQQgBm6lbtFZ9JsmuE3M
MGbKjkR0GZQBjNTq4DVIa3sj2Ji1p5TwKL0F+XcHe7GIL7ArNud62v/wUkg4/KnI
aOBInG5l3Y3O1blG1UFoyNLsBuNYamil0q1pOKHUw3Au4/aFJgfszU/WmR3nRDrK
VXHATugvNuYpVeV8Lt9u1xpk5exKJM4DZduY5TaTTF80HqJ3fMpby+ea1fnM+Z3Q
vMEf1zeVxY8pxKNHQ74Squ5Uba6WTnBPVr5QeO02rPvhnwaVTbzhFEtLLG0x3PB2
P5fkUGZbXwTY6Mb2FTxigoBtv+VMZ7tT9Y8WvN68iG9VBCZv7OJLsld3tLOHlw96
Tnyfqu1ZJhm5uus2AylbNwMt4U190KATdGmWyTnZY1TA7swY/u+zE6AQ7z/78ApU
IhvpWNdLhEFibb8K4Ctq+SRXXzKe5T6jBo54z8y2sUdM6G24ZMPjVyOk/prNi7xY
+cBTJob7QUEDPPgdaavJc8fMf7V3OkAIF0rmfQgqvvZkJZ1oJ5aEhA3+HEv11g+W
NG1j8Rj8bjmYJnN0qesNSeQGSl0heaXWM68EHq4heTGUnRWU7z6SDTiYd4VRRgcl
RTQ/DTOlWFPF5OtJ5mZxjW1KPmPnAUb4+hz/5BHGb5u+UdizlE8CCcwPeA3y1XTS
F293aX99xcwKuG9wlfmOrBwqiaZPiHACNzfcg3hqdA4AkBVXMZdFttlvVNyZeSQT
kBa2Hpq+LMMJ4eon9Nv3HSxR9TiRpMt3opYLt7TDQO6HLrn0pAun7Lk8OsR9oUyG
P9CQ8apQsDND0zR38KLxXtYq55RzBO5q/W92z8AEm4rVglf6VRmHuZbDv9Z8NE4T
WP6QF7uxuHuygkOUA6xdLd3jp2lpkUV0VZAEmplNji+Ulyq50E73b8VoY9dPVLHo
eDqwKXZ1oxl7+SFnWMNjNu/wGRAb3P1dDqN9aHQLVIOM1XW2qkntpAtkSeuC3i/P
L6/3S469vnIva7ymh/70kWuzdDM8hpG4kcPLAR422qXUgiZPpmn+NEEbznOpGZNW
23GYAh1B4kbzIz0PJYRQypPnGax0jy3l71ZMlLzZiW0zwfdjHzbzSs3N8h1saQCd
9WUoqM3pzaWRi/Eq4kPQUg2PhBkjVFZCS6KgBNOoJzVtUDTsRbJGEcmyC6kTfNs/
merzX3ENlILVPb5BdvPajcTsi7cHzJfTTtm6eAJ2uM5AX0E43dx79n5sGVnp4cDl
qDd5mFw+gBKd+FiCQPVsdAnPmQ2HngsK/+h73DWLZHS3XhkVz7O3FfSooO8nTjlv
NvYX00TrZhhUvU2JPkJ2RuDVZnItYwqU0Sl5xzUUgbfetjb2fRnNW0YcLOSPYgXL
w0JcIlD9W5gjj5vhfEXYiQMl0cMvkdlanuHN4T3VNt72JdSy5DLkzyacRyECHreP
Z0xn3ZrRxV0UK24lY9HgTxZ8tCyam1Qzp2CEl4/yIgt0g3ppd/m4rUVi74IrN+5K
QkctfMRyGCUvrc7ZwlnQbsmHkOeP+jOmqdOQ6mMot/z1x1dnolb48mCQWRv6Z2OP
75BwWiA3ZvuhwU/+9vQFkivUcaTe2vAlzIi1V+qT/sGWTTqS+kwxZdrKgPiWTMCn
xJn38aHTbuAV2IdeC/NVJXDqUPbHVlTa8GJv2kuX5wFNmD0cliXssv8L82qgHbs8
rT9FWPhqROm8OMpOOe7i0kbg62a42iGmQmdXviUMRRP0r3bT+hFJWJ4Xo6KOeC/Z
BSZfEjSUUEKtcAnCJs1I6pTI3Aruv2w/iBuj9C0kekjisbsuivgjIJdR52rNV+Zr
jPckKO9Z0n1s+ocxkXRr5yU4l/bHRJFTUG/57u49Xc9/1kSNzh4EkO6LrQtOrZxK
fNzwRjw2gdnElcFrif1+igXZGm9B7CGcLctZu81M+jGURdOzjXJ3Fec2rfGPd8OQ
Os6fSOTkOwiJCnjsQhCc8Rdwpepa1D8pGj8ZNAu6V/84XaOuQQjgUSof72PfNkza
mI9HvNvHM3V6ZziQEp0iVLObTIGAZkSogTn+kIXJ5osM90vG+sepritKsEaQAwvb
vcD9Udg7Lw0g0BsyVFPoblrUlY2G2nY6sGxS7ooPqgUU1putTRnDX7xBy53YCKmN
rEsCJSGOb6L6K/6GBG1AIbwQm5KSoZ3K7pBxH449/GpLuOlJGtXMtbCkBJc5l5I5
/p5q8Sbs0tklpiX5A2GLdVjuh2joIZENa7GtZdm0IsAZ+4IYrsn8waJI68ZeLGi0
9XbBcZ4MrueHNXD9sOUJXvhHpu2EbrvfZd1uGhmyv7dorxPLg81iCU9O6iBMmD4D
6re8dTL5gmA/YhAqfjpk3SL4kBpLphF58Cm3NiJKPjhtqVpF/9Or96rgND7mEwos
B0UVnC/XTqB8FA54XutN7TDaCHFQZE/eOeKhrCavVJ5ZrOTlG+Mr0DGtz7lRf0mz
981vMCL2RShsw1rarqjomKWtOFbjaxRc4vUgDdtHR1kyYWz1h+6QefktbcvT18Wc
eNVBQL3QtmfInh5Gk8SBjYQlUJThu1QHnz1hQkaq+PjN5ConoSBh2DOPr1oOWB1+
MZxZnkhlO6bxBG9mrZYhT0/98em5hNjsHExQLdRNvewae8QcRNjuNFHNlsm1E01Z
0nhkytv5l/oiVAhkqhMP83Lq632V9K8JnFVvqEp5+MtdadK/TsUDSEjbdAMm7oHm
7Il5KnauJPBz9QGuQacuN0sZcgHoMi6qrYYt3yIa3519V2qArdnYIkkO230p6MoP
krWeW8HkjIJo1tw6+2vwm/4qTu372Gywy932aix8uGn6N+3sltZLxIBtso9MjhML
QC56CiyW/pUPtuLHDUzGTSscy6jpy+nG8IK7wKDLcGBX9JtQFMGIL+T2+ltGX/fm
4PadZod9guAXoyceJddGkvYluFfHCDKWrCUemD8MYol072iJeQG68JeRKkWfKS+7
zkvmlX8LpIv74h/l1+dqegWIAAWIF9rP6jagyyfZ4Qs97d71odCUAZyOWtmJ0ZP9
QatVZikpTaESjfscEyagA8pMsQd0ZTPT5HCUsQkLgLo1wtU6xL6v/4sGXpwMqfFK
EzOQkb/WrXVYT9vTVuPvonzWwC+V9yrOXlV47kw61G4vExGITLfWVVLnqb4ZlWJq
gXL+KCP3JbJD1MVn/Z6ZDcp3I37UC7gIVWmd4HAFtZwzfDrQaVMDfMrzE67r5MSV
PDYovPbKe1HTKeu5VlJSFfi2nFiX3lJB7FTLf3ctuTkXF7iiLQeI07QfNTq+Hetr
tF7yFMrcXFaMrRg/xzRqlAX8nBPtOLgZATrnkDFWgEOxHln2+0lUw7Pzzam/Ut2N
wtA2akMC5FDpGg+4DmM2J28SYk+WAS9BOm4D4ff0EHmWuPIENqN+iDFiFlx/n/lp
rO6/6wS8Y/fqxOrOxz4OXa5A+oBv/5pPaLaqHBXVhKXmtIqCSxLsFDyhOvOspO/W
wAcSmkazXXeyb94PV77FoPKc5+EE0yWzqy4o6g75Dlc7InbfgwovJ9YR1Gx79TjU
gj8itqrzXIRwpYUiWmKaNWLyI6pgZzMsGTHZwR+ytkRv2DpbXqx11g4ONKXgAlxP
KwVE1xT3+5OfoASPk7EC9QPfLTpXQ22Asz3mI47Ww4TKRtwLALgXUnRCfkJiniHx
8oTP452zvxtJlWcs4/eYbijhF1sPWG3PRlKBsKzE9+ZNLpvmRdPsEy6DOwF1Hjjm
sovO76H/eDKvCZ1awImviCY18NypIvXL4qztFq6aVCdEfVW/RatslbNp7zTgyv2a
OTMTeMlPju8WZzj8Fw+tD5J3igYC1YgbC8NaMB9Hj3shBvFwj0orPf8uU3UZuMYq
ePZUwMhu2d7w++6kBdcV8N0JvQ1/S5fdF+noE3GAGUeQQhXzq2rDDwVTSIKFM6MK
Cjz4V0xnoi99K9j37x6YaFjQWDiOY7YNggE6GbQK1KPY5PlSGE4Z6L1IK0xkK5gA
TTWiDtDtHhzgEK9CinNhp6D7BpmxexD3yVcGaqRfjx8viKi6WipkS7XGD0ETGBT+
MFRQOvgBoxSFHbGIy746ckoLz61cG8B3nCiLChdjm+TaulJcuhnj9jkboKlD4iup
IeH06/X+lkm1U5pTa57+H2kpbraBSbaHfbg7jFmoZ3PJGAtVlKkMFBYeQL7PWAK5
ECP9SA+74CLpM66xvhQhh6inleesubx95N0GCiQELgE6WbIjiPfZp100oZ2GlFTi
y1MdZd0XcW4I/BiRUKWAimomfynMwin08fj6aulBElV0iAnKojuA0cMzxTiAHU5I
0vQV+UB9GH/T3/NQDnNguONYJt4uZ7bKKvGshLYoxpA/ssJyxbILuVLadRbj/VVa
KAXC+uh3e7Ub768kcDymOnTEFa7sz1HZpL8UGdvf7JnBeFrMezlK3/sc414SJPsq
ixdCeYoxM2zVBiIqRIgTMDXD/53hdHo70fQNtBDgRN1XfgUKpxTF7eE7inD+ymID
q6yCfdsIDfUXlPePeWAz1oqgI37pKeYTWqVS4umExoCG6xDCxKaNix8+fzUBZEda
FSYzYijsZviIpsJl5ax1FNGh+6CewzkmtaTAnwxkxGiw4gOt3YdI3Q5Jgetb1IEB
2oxU0VcMSFpgtiN6wbEpxKLfK27Qisy78qAj/VTls0Awv+G51yQNFna/STak3+9p
QgMX70U5WiOrBw3OGMHZGp8T+8o6+ZtRtgfUISfjqK0whjPmYEM9716oSlxKTeJD
p9chYW/COL6wjqsBljkOALMcEPu8gPFgieLKbXIkEoGrjUF2bIlRvLJAcd8onIMF
hmbnEI55vFtpOhlje6iHT0eMHKPG0WLMG7pDcJLEe7ccO41dV1q+K8aBsGNLOrNU
68RQJ6NkXgZxUSme3xSD0nBmfY+O/pWcxpOFZef89SW1wO+axY7JUTs1KGrShMQe
Zq699lJGapQkI9DYSDm9OhFhnyRWzUsi5Kq0FK/nt4G2/F/6xwGr2fErLiG4a48t
hOO4ivit9YExnN5gSwnkcjUo5Zxv3hH8wl7mkOFFw2zHe7DnzxRdAVfE/WK+oXOq
Nz8kSw3HrElTzIzMdHF4ksc0jR0ZqZZ6wH+Pj6HyQXkqZaIH9rz23bWjFzbzxgWW
3p+KvAuehkQMisagM+SKNd2R6WkFc4FwgXwzhBD9gu1LaqrTx7jWjjg9ooC60DeM
2NytLRUdGQNdSBqES1VDxKUK6gwgwf7jR2TEczX/+s/MUlnjJ2Xl3hUDerWWySRY
872yqDEiwHbYXJqd3tXE1pEd4bUtrEjhB4YxIHKELUOiN9rMDFT5w2CdVI625mTB
Tc8rsImXmIN9qwnOJjmYjAnEoeDMuK9xj5mO8NWYap/LVfkxvi7vKBwIFpkHuKz/
izHTy86tgYW/nvobnbktiJrLky6sUFKU5uNaIrQlDDrKqD2iak1zdqGpouzMM93/
z2RjVbXd+j6sIqRpz3VLkPfa7B7A9KtT7Dp/kbnaR+hyQ994URvdESGQu/aNoldv
ixioMHQSecPeawcfWFWUdxVjNQxBChy8qa3qViBw8Qpjl1QlQPRvjHUQld2nu3hs
vmzItD6hie5UUj3o498xgH2R+Gb1Tmh1YpDmX4SAXO1gzxhDgKICvudNvlaLNZo0
eVMm89ucsRzJjmMQf2nL1JFbo2rsmlfwnCptGBIAUdyt0xJV6Q4wub88pZ4lmBmu
/0/8GnQMnafPiNWwbkX3hDsnIjn+2o79cjJG4mSG5DIiaWffcp6PGchq3eOyPV13
3FvPY5Faq1gIasU+Fx7upVAA0MxCV5jjyYrUCiXWLWAY6csLAeBO5l4kUcZsbl6m
s1YGjL3+hmXdBlSt1y8cYkcG5csbEkqGFbmsfGIfMAJOv+R8ujBmAoQjwo++Mcxs
jFmo2UhV2zVFXalQV9YjhX9gnTE05jb86Qffxjlfw5isgnoaQ0e2afYWttzku4ZE
WQjQyPT9mMt3CCQR4JgV9IH3nfNE+z+CyYUmTCqc0LoQmKViZM031Zg0akid+MIm
98xBjj9hkYkv9cigesBIUhxYWrwYS+0RWFO6R9sBtSEJMoCKSES6yZRZrKZ7ETFv
fo4WqjwMcnrKcYvjNTcggasQzBG45JNh6k7iP29VuPGDCYIcMiSD7cOXuKG3U8ao
rrF/sTV1KJ3sMqSsayUnkrYkYbAe5nZvcWX3EULGwsEG67EtxZt1riv/9p65L4C+
EzxqZxXs5fnVG+aBEqJ4vbK/2jDinqw0VwP/SCawbdz66DkoaGg6v1ztrnNfYjij
daemPH4cddhudLWs55my6DVecxj2n14bZ19shg2SjOO0WQQt3+WtiOMiLHmlytu3
zLyaSwm3RhjQuM/XrbE54O2AOhRt7hXof34FoFOI4Bi/lJCBNMHogodiK8/xtqBr
wObPQv/fw/nYecDGEwi8FUWVOlqZczKjiYNesouWwJTIVyzKOCTLggJO1ssv/OwL
OaBosWyhET0hW/RkriBpYo0OqFsnCqLu1xnvsd9UsInTMirgRm8oTn1nGpq3/j9v
CfvOhrz/NZOnclvbZXRVN/tB5/R8T9ZxkB8SA3wzDsD4jM5hPSfd0Q/blBhqZfxa
9R5Jjq/5o/IjBdafiwVvPlBANZp8z+5UGzyHaqVrEAPkOlHeHi9gkZItKfqWb4+N
e+Y5XRvbCWZsqCPfJIAeH3wdmqFSlUqJVybXSEABWUdJXmOyUooVGH03LybpTfG6
CCUEJQ8Lsk2yaQIqt0Yu7h3Ox4dJes/mexgerwyWDslEq9kar60cf5QGGc2pmpbs
jHnG8YS6RkL39FgNlcu9B2GPnQjePrfUVmeLnwxkszdJTjpZllaCr9ZL1SoR/ov+
yy+9U+A60yQfcEtVuiim+GbC07BBmOXPJvYACXJxFluxy2l2Qj++GIAupYiM+wF+
mGhbM9PrXAbxy8ftXAgY6jjgCXZc70sA4rTnYcXGJpEknwA/pqk03c1C4cZjxjkR
Xihv72sZbvt5ok8206R1X0UP9u3BhEDdsKZnPf03ozHmZGd9bLsgk5JvD3LaCQ4e
eWOzwNJiymqmq94DKlp2i8Q86SmrZgIDkzk+xANH8N7yLWTbwMVIlh34wx+ZglBc
f316PLs5YHh4oNmJOzUMbbPr/d/ZAPS6cwNIvAICcI4HxzkKZoKVzFVE7ji+yi0Y
1cPlXwNWC8GVE3ONmuqtzmBv61Q+k/j9sHnIuZa2n8/usGc4pbV0YCofioOzVv/G
VbvSiChm8GoIZzUJNJdb91cIrYnuhLOdPEcojnc7M2YULdzwDG91IKxVbn7MJkPt
BeWNCLTvjYNLL6XjQ2WrNpzlO3uhGhUi6oKEciEl86oLXfIJXspxUKY5Qphx03Gu
x7yQk8yPzuTIqfvegcLNGUXoI1nkufhJ6rRbBVLtiLx9j29Z+bG5OCOiTYG5+5n6
FjQW+ZyS8ozSGYljP0osZJnJjWanBzhe5jd3Wpn1hbEBJoIaPXczCLFjNCqzKB2z
rFNo+JQBnYnigo29gSY27EwVjl3jIcMQWGlVlNCFnyZGJoceZQ6cJb4xwZRLo/85
QfpQGgR3ojr6JWQcpQ8uaEYt1Wo9GeErGysEI8E500zKyFXeI+ChHC/yw0pT4UH9
xApskbCx6PShDNdi1HqjWH635Te/jjzpK/3dvJnxiFcTSFdQXSsoMhysg52Y1+IH
hqEE4s14SEiuVhohAZLkqhUJhGrkve4NRSHlJrU8RMPX3tKkOhunAi6KvtltL+cj
HAFsyjWDaFm0Sow8r70RG6vPRgXDjK3HPbn+vnRU/rXhVvJmpYBBGbjO34LEXKXI
FLgwJB9bCYZHfEziotwWZKtfV2OJiOuWCZ1/cLdDkAZfSS7TdmxqZFtytk+x3tZX
T0G9FYYogDahu/2zugvnfTWdjWCTCDeRwUr5SEWvb1T2H5B4QzuoF11a9TG6hYqt
77KgTxaWzqEqfpVabhbR0W/dNhr1qB9HnnKuTrDtT6RcNG9evewDbhMW4vH8YBVM
8gb8LMDSojkUJneQHcf/BOn+hJM6OkKg9bTMWnihOX1H/ZhvqhqX6XS8N0XKe1pv
x1aXgl3T28iRRdJ8bApnT0l/Y0ycJrGtsXRvwOzfQxKgPWfvVZ75IP7+OpSOnu0o
dhBiRzDDCmAuekgXkxgmxb1ZjfnxiggefMRAhitwjN3Iys8wQeEyCAfLsxalkzTp
zFGgzcMO3uscvy2E1L/YXVL6czwEsgFcHtzB/g1qv4XuVeHnCKcgXL2F1Z0e0iu4
SHqP3+2X28daPNjSl31zdWGFhcQzyWGPKKHtTfL1Fi8SKdMIgTdufwC3Hq60muyf
v0mCcWNxHgkEFVTJ8V4cOesCKD3awYzuyGWWjfRiuKWPfg2oMGFLe9ZyENjeh2TB
CHbklOHd2xXA3pcw8uCgh+clornNZF9qQcuKgjwXNJXGXaNCpmXCErbUkXtJ6UuQ
YMyaxDLhFlhfjLyPlQrUJS3FvC70wHVMRHO7aKB8evn+qunWB2h5g57bAb3KJ1e2
X4R0XvlFdnc6R2df3L7XXUtvR+/Ae77Kgrz6PQFSG25t0oEBbdz3v3XwwHthI7LW
3wZASXSn6MBUaTLac+JMmyjeMFOfU2iDLu5UPPgFcREgCxYA280EttXKIvdvJdML
4dfTwNDKSsnhcoeG1tc6EPeii652QSzyG9eqVm5So3fPrO6qTyVTapeZ/b6Z5vFY
7LGYZNpie64v48I0O78nzA8hOAG2tqZdWWj7gYCaOtI4H0o6QXwDHfwxoXWNy9e2
+NRC2gXf569mQZ1ecKiGqAm9yamc0L+oFkVY9N0NYkxsZQJ0Zb+07DsdBzhOL2SW
7FcWpmwhLZtXwHhh6Yh/BuxN7fZpKbmcYx4E0FU60NtlCYQ9bdwW4rbuKT8DHDI1
RFQkzNG1fLKxAgm8VvnP7nICvT7kLs4CsIkHBG7TAdHPdXUtVBgYcXd87C4gXa8s
oQPxwbWEi8VbfuOZoEXloLun2+5vV5q+9xzb1UjvZOWSj5Y+iYjp8tFaPgSbNw0Y
zaZUg1AGMhEKY9MiWWCWMk9EMh38Z1Uq78/nueZbBakVjsOi7Osl8kTUGmxcSWEE
onGHBl4xKJ6LgCttoz5btlJfo1uF1qcn6pnUxl+C/HUB5C+lHota8g+ZwKTvYMQc
1ZPsKWBxTgrJ6EwgNAGkBimp1j15Zu1lRBZZEV+j4yiGnYYISQQ2O4m2vPr2VzBo
aTR4asr3HAUvV6T1S1q+XSo2hMTIrXx2n1tReRpGuxHiCc8649l+QJ1osHvd5MGj
mwulYOUpAaCc4q74v0QRxrHbs6LIyeD5Neo2ODm7RANLgFp1izD9WsNrjO7vHPiM
5lItY3WU+9HNak/g+042FMVkv5kVhZmQxB2HuWu0jy6DwQi0HxMl4OVCfA7rclUJ
PZMLjZHHk9RaOUcdyCdTPaiP5woM5YY6Anqh0ntxnn0vZNznjk+VHw9Y+GjBHHTT
CBlUE6h4HeVRTPmGAcnf9G879gv5D6PXHOuGK/g70SsZ91ZTFls75et4rsoYDybc
saIxqjPOBgJwXuj3V3fB6npY+r7Dpqy6bmtV5b5ET/RR3ZqwoZtXY9k+PZ35tOae
2svzLTDFjAXLdgMc1/2PDnY1kJyu7SCcZvNVAn0wL5C1StxV1s6E89xrq1CmPOiF
UONIZ+tokf/K6B6FYkU9yO4d3lJuzw9GacXVsd7DZk0xnxn3wbfsyuidgy9pPWK2
gEB8vlm3OLbtdJFgorRKJ8F7yg4LGz0n6J3fKCdHc/Y3IvJX20OZl/maVTSsZyoW
f+HI+Zllrov5HnqhGFUldFlqy5AHLJ49jETKKyJBA16+JnLrsXQXS/6qGBcL8wbJ
CVCiDUu2DTxih+xYkwz0x4KnpYBxNrj5n4y6kyBFjKd5vr9d1lgxaNADNRz4rGRM
izS+wfCtQgxmchQ/daOvZsf55Y1g1ILFG2D9yV7dQiE9sDCmma0SzrIGIUcoicmA
QOlh7/CrC0cbQKTJInnVI6PjocZY23788mQB3yncGFjFT2bzQHnd45Z3h9BAWCNn
avyeeSZp1YsxQDNje0/X4aQl/UrsxDyzwjpZw5QaKaIb272LdMLSO12LKSe/lcxw
3TwVYV2JUVC9jsR9iSNu2GV1zp8yHpgGLgOXiaw+HvdX6vLjWXkeIWaLUnnOWkl4
Xbk4Ff9BeEdB+GrPYZBOuMCSxKvWidLoIOnDvAuFzseFmlS3NiOk8/Dz0FBo4axA
KVlONb1/3+EIfPk5aKBoxc6TFQFrEhYxlZcpDhODJXwIjZelLTtHkOjRdQD+B1tX
jypd76zZH9GhN5mdL4Ib/aPf0b0s/JgdAo1LRt2RaN7Y27ehwGcbgtlAZfkAyiO+
TsK2Kj7IZXF7tFJkggN3ZyAAXqptISQITrpHpphpz0ZPpOfdgEZ5RbbGcmrtFZlr
jS1yjYh8LiPunGhCTHT44joCo0lbOVY9r4uQad5XW0AsquZk+yjtlnQ7/2sjKcT5
MHtvDsZTCB1ivpxtYHmRGosby6k/4RMzxY4GWlJz+EaptNIIMiicFzNKn7DYBEb4
AqiUmCO2maW6aVSDA1AL8Vbgr82QTI81wjHkW6yZFDJr6fSaI3l9URBwjA/Pg4e7
x/efMtKQ16++77/4Hj4qw1PhphCnUWGZ3vOtIEiTa94Kce2s2N0YIe5X+KldctDB
5GuqCJHUpFB37k+2a6zuS5dK0LjNhNMq6fViWVNmatcjBBEPiBrRXP7RyM3OIsnM
9ZIWb2ISEJXoR9+JrurUTFnxJzwmF2Xo786kfwt86zsU+2Kj1hjmt5HYRCNbA6Bb
PDZwjRqMhpwR/S8n8Mnnt/JdHLt9qs+v3Ihhz0pgKHRTuT/o84THarzCqv9RLa0f
OmVr39V6BHbqHQN2qBpustxLzIG3qCrBFRBxlsTmv5m7yNNHhhELByyzzaaXtXd+
RHCTniyPwMLcDIkz6/XkM9eYitpT7pwBACXevGuRres1VBtiuvCbvTDyAfI2vudV
Lcw3AsARnsSVkhlIpEn/PQ+5BBt+sqhQYuxzHu9dqH3cOsKl8LIDZnsW76fBWzO+
krZgAgimC6GxpH/y+uLLgoGXSBfDxu1M5se4jIZ3rugtqAz73KHMpRWdvDCc9q0g
29GUFdP08PexRMcHUDbL1WGhMpsylnihG0rTx3pTQZI9R6/aTU2l3vwPYjhWO405
lfqvSv8Trg3eVn5sJRoDQbxWgytY+vIX+Flq/y5RV3IwAQN2Akl2b5liysBqSA8w
ocml6P9t3v5YHYtgAE58XE6bCX67w5kkURNk+MXYMOgkCF7a8si6jv5twpg1/lLz
up3AhnydGa0SP6aHYZA30yAItd51oTeYxJQmAcN68RrDXqouoiitzoiz6/4OuZs1
q6e5XyUW2yXZPIVSRGmbAaDhIY/RJcv/KAJjC1O6Kt7ImrQxCBS6f50W/NyQxT4y
8280qwLcLdMzU7pufK7wIbipMNPGSeh/0gAgVeZPbfTcS0w9549GabDiLew84fo2
XUIFlRs1MANyUs8K8lo2NnDKAzUDSI+K577Ud1AMf8TNSzQ7g/1OakoTHyqiXUBy
u1N9DgOS2IIU2C+1VzrsFk1B7jX/Cx9PiUYf2WWP/Pbim6u2rFILbYQNIFcUMgsx
YkM1nTjaEV+miuZbEedd1yFlIVp6fezxW53m62MzmV7YOfREeqMWAJUccPSCl/9p
WN8397W5cVecpu2KZ3hakv6ouD+/Ev3GBiBpXjXp4J4RmX/zZVdEe4Iuitg+wVyW
lRLl+TOY9gBcD4S9lUZrYnwPWljLhMhh9GJk1V+z2V0XQ3lxfdONF5XrGQ+jMYtO
qSNUMpd/V4SzJYVgmSHsoj3uR9VtZIT/2YQ2t5ycDqrq2upwNcXX0nGpyvBR+XIY
RcpzdqgZzDtFLHor1JgWHQI8OFmSDlTA6RSGJO+Uri+XlNn1sucWXng0ziJbaQ/j
6yz9V3FWRGsXM3O9YCvpCMwGDPga+uDz6oBsLVpxpFndUGlWkL7LEM09jO7gRcEw
LM3eeGFkKgZLzY4S2kO1/DINQNKFzlvdEC0jkXu3LZOuuQ24QILGYDhlyviYlOV5
AeBQJfdqMxmherJsdDhEuxJf3qoHNSwp4+hGzTEQERESpeqZYynuYT9y4I5BZmeZ
1aILdRXYY3oFIfc6GwU57rd8H9Ppj67TgQWxPxb2a2CZZqnhz5QgqSIeB4rpqACP
/T2FEg9vW5KXa0dTHJHFS9VcLmSCkXEwHYwSozyBcw/od1RIqHvKQAMS9eyVlcbT
wMqkW4X9lY/M/gVTcKOLWafYRxB6apjZIhnIIodi/+RwSNqZhypuK80EaxiZZkeL
d+aZp16GoccwIPBhcXElNtONJTjen6JkVXWPXhBhz0sWaWQ9RoIrQuy71QY6Q0oQ
dbzM8wW7DC1aje6JqQ68GLX4m8k0xTcWbNSa8Q7JBp1vSwldGaUZnSW/wdqlEZIh
2HlnY/OUmGsaNmhcXxzrtLcP+Oycdfa5smFubocJR69unCegoHQeps/bd4em+56H
Ac70b3gQ3Rj9bVNEVe33rUaOAwDJ4k0/W8hFAhSGFZrYZ5VsgPGPx+6/Vup1c91j
Lxz9CqLzBeYhZV4WvZ2qjD++qLfAgNrAg4eQcEAMrEwe7ugJCHvnedkVIzXtMaw6
ZQ+0Y0h8rdQwrGRfX5jbJJ5pwYOlwIIrapuz4+rICJkJfKF8cYXneBTmScFCmDxp
H/dsfsShK/o95HzSHdqnp2jYfJYAhtW5GrmMcrQhi7oJkl/HWk0UJm+QFcL5wk8D
7XQ9z5WTMDxvRZ/sYfGdPOPkzl1EsOt6o9mJooKrTk28OcYRUz4RfWd+1gskxTzk
+niEhZLtpkxO0yLH3WQFpAQi0OCI2CMXDxs20E01VpCv5TvUPkdOAmK0XkTPjt8z
tdbtcLxAoeXSEVB8Lr2cXKtVa28QVRc5V/NXKCMXcE7+ZDfyR2trzLyfs4Uy1cg4
4YYpQzIq409c0/jq5BrezDU9I2AUyqB1n+KeDNgGs2b7XvfvQ/tNF3T8UWmnieJu
drX9jfjrZa2FtZkS6Yt2oUnHB2/DSarBgWVRM1xakk5nqhBAH5LVEodBmsVpZVz4
Fvxr/57l7y5lY1w314S5L7IzGza4xRRxCrKYMnZhloF8lbxUDGAojPM8PzVrFEpQ
LX8qZbLSteWv/eMZKQA7d/lAwO4Q13wBfi96q6Wscdy51WYhFoDBJNX6mS0Amemq
AV1ap/stSppsyBd7ljFjr9PF2STbnkW9p6xUtwayKw4SjFDU8sEA/OOxPt5vyq9z
+QYK+byp0S3j9WqBn7miLxmxjBQ1MD4Ls2QH0saLVhcdF+vb9Vm59xgMmVCQSmYu
AukyLoHubwXJmqwK6HYbnMsN3q/8yOCXXf2RlBV1owsYo6radjGin4jZfg/xi/e6
z50FRUCtYnhMrchEofQMn8cncd1Hhd3B6guR3XTQrBTV2V8NODHxPmpiUQItdKrG
ZATdRfoA6q5iv/hI2L1GaFCwe1roIEKPa/4i2Je9NnZxToX6InO09AEyYGhJ9ZwW
Zjfx6lN9saLxZ9kaQSrziWnbg+d/KYW0zzXst6qZzmSpakA3ZL2w+ClE+Ki+ArtA
EuFYsE81gdj+fB2fhgLQXmjbsHHH/rtnJENr0Pqnmq192jLKciKnXXL/AqunZK4b
do5T+gQ/9I46P3+P+OglkQkM6qg9e9cu2Ke9h/vc2YvSvKhfvHfQjRfyceCc7oxe
qH5VhkmnLlcJB62jifPaLTTY8mXvQk92QuCft8OQumGeQK5eXAjG7PUBlwmOKCtC
eKTbf17cqoE4nVmR+8PoaeF7xXkLhvZG4C/QxNMIze8r72MTS9L62IuOCUIcPC5A
vbALl8JHyeeoayxERJCIdbpOSQDTfa1ePyj6+b2WLnSDb5JofqFj9Od/Oh7wMPGx
NdkYlPURF0oSIinGu001QluARQI7wEPADrAqhi68pH6bcLv+L1YOx4iu11eaMrHU
A55r7g/obBfGCml52L8ShLZW9FIlFQfFtOnEzv0RA0Jo6iHadIM5tIDRZ6jKbJoH
wXeH1JsaxifAI46YfL8jAyys7VH5b5JTdmGBD9lwGPYRQN0ZvfpD6oPivTm6KiV9
Zol65c/d+uNrCK3yrtC2UbYZfLHZTd+J1ONrNAfkBTKFXXtTpd+6RX9W7DeKEgs9
rgSXQ1wZDpbqs3C2aWYxzwUSdNMCWI/GMaBgr+n/FdYBkdpm0CxzlYA97HAdPHDL
9n8KW/SV6keVB57/6wIRn3iFyyKKo9JYy8ikh2q7xTVAtboklZaONcWOhXZABLI3
NQb+YV6CDWQkf73wBe+q5wXlMrg6U07AouRwGXvasMdmFzFts85D3RUsx2X7LPWL
3gBPE9G8nz9tQoEhr2ZoW3jm1SbQm8lCAaonryXxlj5xEMj2gD2RVHpMLtUYjnx1
w4daTOr3I8GmrMdR/rAMp2y9CMxrHCWESmkOCMrhGR6RNQiTSA68W/eIKTRv44Jb
WXSCCbzWiatmdY+PsTwME85RoCNiwPf7CmcaRRPVUhTCqlFmINqwsystiyXErvzZ
HfjPwJUDWPSmM6okjihBSNDyabZu1E7kd8gL0puBjb/xRgDmwMWMrtPEn4FefzHh
DViDqInMRwmhmpM5s0dHkSt3akoRkuLhhOqPcBIfe4XqVeDf5JIqVuIMvUZ9ycbR
Wt2wo4ynYdipdDpm4DXRf/Yq4bPrGUJU08C87FOtseLstLzkJHlxzfZJFCfYD5Ta
Yddcjnu9+7euDX1y8tLXx90k603eJa03edmE99QfdyTBSWNKs0zzlNCNGfKRjxx7
CEkYTCSWTJcwKfXjagAs7qLFbF70M76yQhSJTEwjOOQkHnqrDzlyKfh2Km8IxTVx
6pO3MBOG9RbV5J800Q+/x+y2RVgZC5aR+2gKSIxVSxOTtNKC/H0kHUg8m75jnU6P
n4D0FM37T/D4LyE/poLGu8+LcC5VS2PhfBvrHdSovWFmsdlGg1lKZQfMfBuisdzy
Ryx1qQ8oa1D44NvPGpNg2mACKGzQ/FFnjEDbGWR1r5BD7ABqBsxm7Xp5Pvhr5PAS
UfryOiVwNyx7qZ0iX21bhm8iwsACnl45FLxxfnh0qNQcntifTbZEKI+NPq3b5lKB
Fswd2xbjhX/VoNp528KvGKJOt/Hr44yeiS190NoOhWo9vCKawrS9MJ9/t86O4G2A
tzqdQm0Ik/5C316DB14+5vYa6sTej9WOSAHk4bz8Ii5VNiw64RCoty1lN8PAHmH2
EsAVuuY0+75IBzhEbvwOpJX2N8FwA7XV3fRNnryEi8ZQzCvbfLgqAa5xbb3+HTAY
eA6izxkJgehXhFlYqkHA29QZJi3yGpIIjjbqzAsNX6ACl1aHoZIgJuh0AnfD/TTF
ZiSqMtcS4vkYfVxzm06ZhLIWU6Ep5a9TV7XAvySbGhEGLMB2lyqpjrYHjYctlhZb
uSpn8n3tZwPwlmk7i8VpHHlIFvJb+Rw5HiuPChW0doFaaqRNqFwG/+cFBzMCF+Hg
bmAjPLQQ8XHussOCcf1RxTx3W6dfcvcYbG4W/GBjS4b61WGq9drPJYJTnUGHVVhl
V9q+Tet0ShSJNpB1dXwJL/s9RP5soTluyBQL1nOSZKRhbg13WmVFZnrhkE8twOx0
BpvhgKzKPQPiknxZIq9re5o7MKARhe0i2dZi32TitWs6r3mOoN9fAbSR2QZYr9zy
XXmF2gtHQuzFJ2Xymq3qhT+Uqhct9lpG5vsOCV77j7i9aT4paKMJiP7982+1NAnG
l3nM9XEsHcdbra9DY7Y9pWEvLibVAa5+doVD5Q57c8z+TBElhh8fjt+I+W4kvbli
8ZJfm+3/Uir7tryEw/oW3oVKKgHcRW04fssJw/Z+3qpXxMTKReaPrzbqLT5lr+NO
R254ZM1EwqUKKpw2C0uHNjdZHGnLewP2UAMkxj8zJTMXRgY/DwyVUtRoYJyA9RMF
i7U+e/Yym443y1JztUIeH+G+s2FARtg3Bul1CgLRzQUHHJcwsi5fWCkv0c8rExQ2
8KfqJSzxZNjRJjSxA4Yjd5gh1enyqphsMTggxJNAPILPZWh0KH1GziB4HYFoevSH
+1N2Qdegs5ZJW42+FArRZErFvIcKRhDWoyyT/hvHQbXQ9zvRLLwZvuQXzininTvD
eYmyPPu7iEbrREx1AKlYQubfrP2HVCNDQys4NsOyT5G9xdAFadsBD3mZIZyUNRQk
/NuDoLAMI1Uk58bZqSepj24/TmIYA7XMSIJ5i8SRpiiMijR0H6L9/FPfvklERQN+
+Th74AyhVIkVndEZZMTd1JQGRQ1aALuS4zaEu/2oh/t9B/WwqtGwuaHQBSG4lsnf
Y8Thkw62UuOu+EeUUMpEyDu1HnYEAU8dHhZHzOC6cWP87T6OBqJbIANgZ9ULfRT5
x/R49EgwJy7D9IQEWHC1jS+xeAusoeXMcYUV0vE1xLfc60dHW9/u3rddK6NP9gM5
VDPl96BdAVn3VPsSMwolAbGNVGIB53RX63bKnREGt2cH1jSrX8CcMbgPk/K6VrSX
Zq4iDNUH2vy1T7AjgfIqqw47fgXRUjMe+B0Awf+A7kanlmQUR78JSSNhixWpBfAt
28hZjR7iYX2fv9qWLeSlPhYMgfbHDCL3qeB47MJ0uKQZJ17hDi9EinY9sAn6bJOL
gaCTRahNgbRy4Fd79+2yQm5N/PEvVxXHg+yATfcVemaPjpCeZhNjfMvzwh8tseHk
bacoAh73Q2+rLCUReuVjmpLfA8ON/bQvc4g7yOPvOnElZsL31pNq1PqP/3P4p3hD
DepaR+Yj4W3P5nAKqwcx+cwyPyroNcDn8mGS4lvP91DA1ODdSKWMsJTLM+REgXbS
gOjByQg0tZ3zUnYyhVujvT8o9RjQhE6Edc+hj6S/9bZTcvWdCbpSXmWkcwCUVVQS
1bybh+kSHiMEL7H86eDnFGkDlHoXA/NNjg3OLurpm1sEzkU8iY6xzji5/1TY8LTl
NEafoiYRtPs5YBSYHkvlxih6wtwZi3OkzKzXpBAKT5jTxpDrhAkDDKzZKOp7UPwd
Ky2zaPriNu9apiF15tcF1L9cXiwJy2QPWsSi6aXl7DUX47GTGNqj7pADPJcD3Cll
G+/ZC22p4wmlqw5Fqnp/mvt3fbg2O6YfhGZHskh97OFfZRjrpLPEcgtYc4etSZNP
FksUhTvfXNV5kLbuLLT2Gs08/B/9VpdRg4qHMh5LZ8vkLEjqHUt+3aQLA3IxPoCX
2b1jGVL6LgKHOB9QETPi1cGUUTwaTT+cy4N4wUNjcgdMj2sgYqAjiI6zVpceIfNq
kFnR9ixMRn/IQwtOzXDYpNe7ORXOLrwtIsPDXGoeXO01czNLiAKjq2bcSnawqUt5
GIuQA6S9j+5XWUwnN7l+CNTGBQSBxMXx+n1cKGdIuxPvgtHhYhgiWGSnpMCnJGGX
eZ2IiWW6lzXWoiTyMMr41BKEKCKRMCM+YxdJRxhOvr/ju/Fi3dTDSpDvaCukkDYL
dSfC8ZnDaHJWKh+AXA3d7KKQngRiGwrNbX/cTuCiH/KhTWNuiigT+p8AljzjRwDH
s4WvbArxT86BxnvvMpJ56+59J4ATbJCKVlDGFFL9vhYVCRCZuL50U1f6gg5yJlgV
7uoVdPo0+r4GLtExzDD4mskxGIUsfUPKhyx/IO1VsepBPQvHf1qNXtpUzzap1Tel
NdY09x4kyIqwKmEvU9bqh0MhA7Ee1iIG/OzQjtsP9QcF8XpVGBj/HVGQgZPJQpMG
3xvUkphwWig96S3WEwK10JCvnYyhhr3jRZ6emRINdgpA2+c2y2NoyULBRrxC7Ndr
OmyteSAlxMSa+0gdKYpEfafIA32Qf97q0D0JhNKVnwFDKkEjf05Hyz7YuZ3IvAVz
dypMRP5KlPBgmblljOT5VDQjgEw9mlMCBUK9z/wQ/f7qhaeOKmgePKSuZPFxU7Md
ULrUtTr9XES9R9OIMy5iqFt8brJU6f+2BF22YByvj1Sq5dnDSLlBEcx8+v4V/ZZ9
7EfAY938s35+97rFaT0AFpIavU06RhvoZjd+6/VfIXi+uqcID2WsbW+IK89tmvpC
LqjLHr9k2AmFPq7Zn/KF95oT8eG6lxE7+D1lu1ZayzxGtGFj15dpPXfRWynGIFlK
j5atyDA+zmvQz+RGsVA1TD0drbDjD5Q+/tR3dGDO7vBvcH94tM46n134MtMLCqf3
KI3OPnJLxzHc10Zc+GvFEKq/5sr/jGy4Afu+k2WPgMNqRKUC7p8D61aSskwjnPd2
LOET68QSSjPWZCNNJRgi4lhokXtexLs478DkHMmwlz9ECbIIMZHtmUvN2tuFBxqX
Sj8qtQ/UodTbmI3ZGrR7w/rVtuCiGyO4wSzRL3r2s6s9TWPlKXjhshhhH50xyI/b
3AtsOm4i48vXwIazhUsgjIQ/VnD8KSh4ejRKby4QQKpXlGTGt+WUbMuutw1Dzr1T
cFfZ6em1s19k8W0fxTJkWt74SO4DOB4kcNMYciorTmHjR/C53qbpanF2YITT8HVG
loo1MNqvJouiY9/sHv9jn9X0++Jz2tyzsAYlM38WieaBRfYibRh4X52ba3aXz3mL
WLl4JV5Cpsyc4xhu3NcdwMIOREMb982WMQBIqdq5IYyFGIeBbU1vLAbdIj0Q6bR6
xpH7HiZMczAo6R0jaBPyY0DI119Mhc9R4fIOqqhjFz1eH3H9COsRY8AcXnrWOScr
gPEl34Jasq11FQ5LseZq5dgtnuvL0EGMdPSWiZbtWlt5R2qhnH7fi/MBTAqWs6GE
XDOX6YqMDKu7NPSL7gYFHrW9Th4MU+ghizBK+nYhqAVL8CdEjIoj1KVTwjHJW6TP
eqJwn5uy6Wh+hoyUpT1UFuI/d/EeWJDoTynwGKZ0CKsB0TgHMruMTYBAPIyErvcb
tqeCp0fps6VUagCkAmZgAcgYBqTFdQAiBfLOo1QTv+grXBZE0rI+kRBWUDLl74wy
BdIlLmO8jLO966Pck1sJ58v3420fYvCHuSYXOgy8V+UkcRxDVGx9iEhTtqmsLMen
7jOR3BcLtHsLA3XY0IreB2tc8i3N3DQoyqjhAgiqk8PDuwOpriy/sCo8yN9XqajQ
zTgaVS7SgKGUwJI1ihbtkmUVn5NNSOvQJ6pVWfwb7kIm5fcLZKT20BMeGPl3NwTI
uCI54CF7Rgrs9Zig66FuPKktd4BZbubjS9eIBLTfgiKMptlZB4bYPfoiBKfkeOJb
wozBcuJk0yLlDDPK0yQzi3baepSMZpgDxAAH24yXv8QdhdB1G+mtr172btSYgHmJ
gL4mbzzMRsw1ob84v/lphv1oKpSNfgVqXY1lh4ZBpJEpm9D3J5LdKIFAsRK1tjFj
iJ685BxpD82e35YqEdrlLPtqohMrFZX+WNE1Qh7Fa0PABmAbBzgD8gTkmaFxmH8e
TuzYo9tvyyPLd+leKDKLkIkNyBlHs33u9Mrdk5pOGeSlLDCbf7nvK6tpt6RGKomr
pjv+8VHw777Y20aYEXTaCpmu82CHjs+DWdeTNcVDZbgndLs+5rbUSRya9Cg/kCut
IkG4LodzONJ5ICkG2cqqRafy6wFXb1iJhQEeg8ksM5Tvyh3XbjMGtwDlvSOB2y9M
ZzHE6Vhg0Bzrtot2WyQzWFFzLTW1hLxx805dL+nJG3fRxEwNkNBf+TI75uwxQS6D
p6HuyfzWRQ+hcAzHSXs82LGsXs8jxDT+Ja9sC/LZhwLB/LWcxRN9emA3/I+U8az7
R7fi6gauyQhT8Inh3uNTYtpLde1XyNNgyu0I7Qr+vnZUCIJhH/8OnTVUaComlNZ3
o9nhhfuAdwoWE0R0CztFMAuuG91p2UU36Ropl/gnptNFcPvjj0G2yFPx71zwF8TQ
Ms5xunrccrI2SUECFV209JBuLXS5qAKYIQVEuEH7EQtQiVA0FV1h9yeaj1nzfAYO
IPpcXM7TbcqkCqdBLlAUtbmORi/+oLD5TleSk/IJfq2kTpFKV0APeHFEpANECgeH
KeJtpV51E1SrNydc2cqOUhFVURUHnoBnchVN/d9u+8AEOA6RSn0jMyrjrWSLvDFB
HOwQp5Bfcu1Xfa1CN6PTZ6uF4ZC5ZQEvD2kZFKXx+D3OkZdi/CfW6awLOSnKQQCk
fAwsjHaGKY2hcZzURIUJCND5HrRxwnIBJ22Cw8PV2Ggk4BvjyIIRQEFKdyFLuEzt
gv0ujgcQhtdGF7gV9DYj4ywgQ9ewHffKtqlkEu1YBaLGrVJ+pL/rc37oU32l6joo
xoAM6qD7SYVr8CtWr/p/zpXYEGyci6uBTFxskOkMOFz3UBQPGbI7EUYC0V3o8gll
65sXWYcHDGF9OLxirBVhgiQBDkJsggdQggYtDDWDLh1DzHtORDU/ZUUZqXMLQZLO
r/P9pM1BiUfjuFRwxcRUUgGjRHdiUADAGI0claGh8GpKLAIIviwyet2hpUh0w5xg
ci3uxZwwcaXf2es0OGaWD90BqCvhVaMl30KBPRJItNryaBd8zT7WBsyJcSIa0XxP
rL3yco+B79wXsWy+qKOnbqXKGJhKxKNIVwN2CUqUA4N0o7lgYHAndP2m/UemB6yO
te4ZIlsKbeYGT14g1eR/4wEucLPUow8S0WbbQ2TlcaUBnU3X3R/REBgoOVZrk71k
iljHS6Ogw8doKxW/o0aSXfw11yYXTW9dWHfD5E3t/oacB31JA6yx2mJe9f7Tj6kS
hes4Ig42WplpUTBQju/lnHmVACDVKyHENPJaC5pDqz3AS3Yn6B7uDaDvcIG8gGXz
qW4ujqj7dUTto+62Cw/qg4wf0JLPeZ5NQVYufeWffr86SnW4lmNh7llAlWW1WCta
G8gaEr9NkiwmXYy6i+ZXsjXg17V5Pq2jfyJ874Lg5dkGRlj3zj7zT1FJmNH0CV8y
gSrnLoQ3BQCNNyzk3Pd41GAyHHOfkuVveUNFDJ54fC2TIErSZYZEIagALuPP0WAI
e5Y5AKfUhlAXfoUJ+dzoXydCJYDofOY6JPBsQQw7PGkdhgOr2ZUBdkgtXP6A9IeN
BMKr5iX6Jbis0S2ajJ+O5MoGk0a5sW85pNwRpdXw92v6GKMAIJqo8bORPLrczHMD
ebK8SzPwzMqbcNvc5FCzcprJJ2Lw6WVK8d0TscQbLADtoSfCSobmDmqgfG9iNru3
7zbmFRvjBFSU9vqZxB7Bv7KSbLWof8gngt02s6v31a7iK9X9A5mncNbBLZVNDPjC
t9j0zAGg2zCqgqbd6wlQxW3nQtuVW1pOahL+mE5NmMoOSa/NLS0Fwg9++ZclADj2
dWRkudXTo64JvBwL++o7vljGzIZ4HQbvXwcwqT/eWO26dkNEy5QZrcIsj5hV2cNm
Rtd4//heEQYqlJeuIQzaoJ5mRzMfNapsTacuml9m36vEG3xYdzwOwnPvixalOP0r
hKmyDjP75uwyGcDQx4Q6Fs/dZBbnsA6MTAdus5I/f1tNuHa/LtviOwRUdRflZDNK
8bppjqcV7HwAq4uAR5qb+0/zFQfGFxWcU5nW/skHA03xSAp1VZjh8bXCIV3E/Q7x
VTb+kwXDjWkwYKbL7fhwK5Zh6giWqWBX23eE81a93p50+vEeLoaq+urZPdNBN5Ik
Cztkid0fS72boRW+kxPlO9CS6pjzafdaF9AQ0NsihC6UBNhUJ1X2X/66/0UyHSGi
5Q4TIYlV2CKvuzUiJxEKhybtHRKBlw3pooYD8E4IAcMRJboGMyehCJEw2GjcWGFy
JLKhdDvLFQi+vifJstuFQ+FTMnuAUbjII8Yhvh1ThSdXmFTtpZziYQ+3F5yPBbOa
LrmeNLpv40URJ3Bvik0YZQB+RhSDKxRH7u87R7NmeQhqTDeRyRYF3BQtM7P/P+gI
DpxcgWHPTNy4DzV/ZkZDFXGMnWmhHpI5EVF08jDowYIsUc77M/iCtUzI+yFakWvz
B0/hHipZVJKq2JCB2qsooAmQyRpY8n4sOoWS2OgToZGogCHoBwY14M5wGoI7sQPl
/1jTS6Mv43OqO7vreZVXueYaZXKx2qu0+HqVrqFuEJxmphSJw2kWPE7VX6nMlk4q
M91upWTHpjwG96jrk0eLhudLP/KrI99bnA1pk0euxpwsyItQtyNFiyqQEeOjiIMv
rgFN1pUFGZiE/gpfh3jN6PcYNk7DRLXKdDBabQupE1rS9XxBGDi2H/qHlp8AAIP6
kkQStm9TR04VC0LhDOU69qC6yG6mip4wvAYsUJSmyu9E/N59hLDvKsWJVsi+6rqA
9ArpSRWgnIX0m6p3jh3QxB1foS97pcQ4XJZ8GNrIxyyIKFWkJ2bHYUNMbshxVpw4
K7d/TS7swOYbJNz72jOWj3UH1xDcOaQAcSuwG2Vb0HLOgHI5A6WIF7hfSa/ydKxx
jL5cFnoGXY9Kg/Z3wcVzZzJBbnIh88liEn4G52yWkg4EvYgrrpaTVzkhg2W48++0
xl57UWw0OS2m81K2yHk7VY+UBglqmrbLH0b6smhYbmlbg+HyY96r/VPNyt/EJJGe
wQwV5vhrHa60NDN46GL6kgT+CjgzgzGkUvOaG313IapYqRbafrE8iy7upjajuMcd
i6KqMkufULn+MyXNl5tgnUvY1SnTd3jF+ETul8bWQjb6qPmb51mKpepQCOZ6Srp7
2C4jVag6Z7QPEfD72AxvRP0Mya4ICGonLGjFKB6d5GKAtSJHNazkPG0wPZn/UBpP
j0TpDUaf2Qk0YODs4iceI2Cs1tGp/hkSl17YY0b+tpF31dd49ZF5Jw3hPBjnyxKb
D2nrGN5oEQNZTl2wDzgon0V1iVZUCXSsWauMUo4gk2yonxbx1M0gdGat9L2d98m8
w6QLyiL3ly/q9PPM4vp95njeB4K6u8BkJn1Ia7xecEdWNE/c6YEHwUDKe5Fh1m/L
C3l2F1ZBhdr+M9syeEHDKX5YGtVSxYbUX7OoCFPoqB+/pg8PCwpNqC256WEZxZzh
7lLGqfyD0BA/9br8iCVS7gOAvNn8nLhv4qQpYS/8OMIeSvGLBxJQ17G1ZDl0ipOj
jREWuc/Avmr3rPVVy3BdthsaAbwKKcQwj/sKgIqmkhn/grniLpKgoce+rTQmAkgl
m9MgHzwNA7mJIZYYZWH9zizzRL+xfBZ9WaI1MXKGioWfDKaaWtuN27HQ+RdTJEjp
cZttKXn5tfDB0ZhVPgD4DcmgzxLCmP6++ttGo0wjc1FYDLRSxAt1lwuHOIPBh5nQ
5bZTwcfhrxTlSoPVA+m7+u4GRh1JPqiDRkMzjy/opGuSC8yAfGb2I8RTXx7fybgU
njNbhqvLZW2MSonWC61VMtWgqYhHRGqNApmAy6nowAJSNDsqsJ99eUNaCBXPkBwF
DgBS+/nALQbObu0OPYQ+klkFcgGfe6zyV9DEpZVlPC/bGwtLJ4rjoFok1zchChbB
3EA8Jv/6XIRSanag/X9nzPpGdnLgSJaJXyiaIsehiX/mvD1GzQXvlxH/a/hHaJk5
8FIS6uEkQx2V95ODMH1hwuLyfaHTrpRuVfbN3TWzImeffDH2W5iy6ESTqBkKQNJb
d86PiLkqc8LYjXvdbQDVOt5G6Olk/Bd170c0sSvvcjy00KKg7pTSwgr9mP3M3W1r
w3RZuR8+FtFe5VikGUspyBY1VbMwazwRBEdvJ3MX92cxqcn7GemGf+87EICUBFn7
cxCtRXjJkcawv6e0JnSFe5KakK/KViwfxsMXoVfGzTr+kA9sbXCdDMHYLMnVjhuR
lBj0NuS4Mfnwv/dzoGl+FZ/WgmT9COexU+m+/ehfD39xVPQ9hvLjPtsWhAyIfcrS
ahklcZYAfdAMvTQs7pvXvDefh8VI1yXsuXJOG7+jtvBKIW0xV9ltjNgSIlaQGWpN
xMTkD6tstEkcZbZeTvS0QNHNKpurIaz4sjBEjl4WS4Ua2KPXfZmRBwVxXoOJFudA
VgB5qLPmosChH2Koh5IftFJeDfm9E5r08KZjsndO3sw+ENnsC4NLd3khOT4fdsiG
IKjppUK+VndiWFzV1uVvQp23PJUGhom7m/YL6Z12+Jt8WLfIJO0bbnWNn4n0xrNU
vqqD0WNlOp/dal1/qrg/Vfk15w7fAoctH3zrUHO+FUM5/H5onHKws80JWmHfqKSO
qQjd5MrzMvgjemukeGDVrG3S8WheLpWPVTzHSkjDDwzA5DdPcwRDYJAPzvpnUwMa
UZK7wyDaVLmW/qRiMJ65qN848ijOEeCwbmINjrlnakJpXJvifust1h262fPtqI0C
Hr4XI+B/ER/sUn+m1ZnzBih7J41EmBfy69p7yjzxo02NRWIu4/JfssbMPV54TYW/
tn3L6iy4yXMBL160ucc4xFa85gjXw4kLCFU/S1if2aCKmoNZ0ZoGI8mdfH+ug6dz
SlxCXnUVju+gBBHL3EJU01YqLL1M+VsUg93eDbQ+DTVbCAcqpQxotJej774wkFPo
lmdFlaBW90YeoLd7OOrgAUFJMws3ZqFABb0xwZAktgpx4Dnjsf+nU5afu+2/Q+s9
GQyQEeNLyunOd9t1VV6fsYEupFwE00osNSHy6nT+Sbe44jwL3ju3alzB961lvAY2
yK0aoVs2zzJPNdxCUhcJYhYm44C5+pSeCMz9laCl3R9hBBcLlXJum3vCdXLoBH3R
qJesGLzU/0K2H2qegFaxMG9jUQdyfVSRC+cFYkf5/4Jk5HZVFRMAo8vg46blI8Qj
/yj5nqiGoeSPNkLCHZizRdqBtmqgYTVPwKn8QAjZp7vacay4TIm0GTvMXaMD0wuW
SR3V8YtV4AF8cWHO4y4f5R+2n4mFvj1XD4NbLJms87TinXRh8gcllWxkb950wm7P
hoTq3OI9JJTtk2ECBa2YK7wkubiJX8Rk+0YZ/rDCZAAzqR9MQCxAV395NIqV03zW
4HJCDEsDq2JYeOLRZJWidjbil6jJKSJdXNM3DHcqW3cK691IqP4EaCcTx+bDLSmQ
A71njcgoFTQ8W7U1HP9NvAbJXXQoJ7GSreoITLqv1xajrxKoz1kUHMtBnTEqxxwK
B3KgSzfKjUtLTeZwr0XzYzTU0xRdT+UnBwjLMFshJxGLcxTpkhd6O9HF/ZzzqVU0
5tOVYO8INROLKn727iJFlsDlcbw7gefWK6jTfossH2My+md98t022JRVL0XVZXKY
9V0agHjMuBbx5M2Nhc2AsemOgYJhuXUTuWDCxrWbyVVw91mWG7/y6LJ3qpsXwogY
kB0P9Wy2iW+T9i60VDiqTCm/lQQm+uHsYn/jHH89SE8/7bSLz9V8IGbMOEMr20Bk
Gvg6CgZWbzSQT0LkMLpg93tHZOXmB/DF73+4PepUA+ZBOk1+4Q8f9cJXcI9aZUAj
ucnDGqYk9IaJ9werJ2foRo7QnaJJ4pFQ6NkZJuFdxu3VKYohRCe+Y4iAkbvx04pf
LDhh7LMaqoWCi8fXM6F4b31iKGaSaLi79Y7CWoSPtpfQkx8g51iC7mlzAWuRusFY
/pIWqGl9lK2b6w7xk4RFGyBp4QkOf0/mddGCm2B59QREMa7wHngIGI418o92c25j
PkgaPecGwIH/KWsy9a6mDmp517ETj9ySJncErw9cFKIL/4FiTu6ffxxvbPg9MCI7
gkNQ9Y3WvssO0NfgzD2VuJdwWkOvbmQXMOe3T15+BnZiFoPok46iqli/yAcySaR7
KZljMrQ/XnVEQyoOlocMee9IzHtZcT41IXoMwAHCnr0yvAvthtl7kMzEcT8E7rs5
CJh5/858Y6FU0HLXEgp2Y5RmkWX7xeYWUbClalLS2MAghiPIyEV57TcKbH8Ygo5H
jb91b2QXKhnyAwOV3qG8/7UV8cwbKiUJJ3js+le03nVu8s+LK32TuggXBeeKU/Mz
jYaacYqiJiS7czEORdGdKhhkK2MydGT6n1t/LGCYk4KqG4tda6M0AnEatF14wJVs
oB4UTpLkqZatR14s5+r5MPGryZkIYkn5nbJPizxUyXKxMqPeMxv6ytlDd/xvWGEV
WGIRnos32tc5O+6pl7pHlZrEAbt5HD1g1SB1X4Gaiu4m042mhBLJ3QRleoOz1KHe
qYfQl/56cu1TAbSV1urvfUJ1VPMqeL2X0xj/gBVS9QHOCp58YQjCbdRhxloNLaOd
cYeTv3Y5h4+mnxUWArXRuMP5aH7UrLbxv+RNKSF3pC9UY8tHNBszi+nFqLBjO955
NZ3D1WYb1oZPOMAVXq65VNA/UjnW/9gGBUBg0FueVe6KaVlMxLnyk9Z+Q9aklOLb
M8GyfnSn/hcB53nWzJvaIXQ7zQsAfGvyIuHvFM6ApTlkhhJ90d5zNiiNAl9as/Yp
CKsANQGbfFHqB85jo7yRyytOrao+vFzrc+LkN6dI9UNPhCyBBuJoCfMZ/1KOBiSB
MvPCZP0CQFiz7u88GlNOSyw0mDWix6OdfCtUtro+IPvdOC83BK9pSWAKTq14UFiD
mR0meVxdpS9iYuPRclJhZQUdXxU2L2ukNDmZ9ppnIlUF/5XL8ME1/yOzSNjW8YET
lFGJW1FJle1h/frJi5WxpgP6MJdech60ViQbq114FA49D1pvdKL0oTQ8OFfJwv7L
lufWsgTMi19x7aN2COwr2VXSgtr59L3HljZ15tbO2+ivIiBAQ6qc7nkfkONZdzLV
qMVruy55O4dCxE3BEebLFhxZ+1tiKYk7MKdAknsr9VzGnfJdegMW0bpiuFBZU7tW
3YcZhZUj2xRnitOIvPJV5hU9KLSlIbaJGc44zF4efqj+sCefi3Df9ab8y101o5Ff
sqi/8zmW7JpGnq3kziX3t3FQEQuYvdYrruRZNOzZXpekRI1W/oaX7Q7xepOEb8vH
OvGl8kLouKjyTBkun+AWaWl2oKyBBucW41SQz/SXa0F0wTufGqOhS1HCAwufsZI4
Bc0aCN3AhTKdBBcMdS4LbWeiiibzd5VBncFO8lzOgHbpw7JToQmTMR12iPiIid+8
UFtBh+jZ3QwsNdW/tZaLkZzQC7/s/UWBEmmLVk6RT8nIIMha0qyJA1WRuv/CbBco
jO+laaoeN5KG8nW7bq+CxItYqNcactAo0vSiMxyDOkSN9dRFmw9r+87yc/TXSa2c
HbMtQ4+GA4aQPD0ZNJ9dXeiW9pWrrUMWoOqqiuwoB6KVfMO0SyKrw0IInfaQWvTD
ApfIB6kii0Dtylu7eHa2d2LDIXGcTmrfxMK/wX6zeB/Y8Y9mpdiEVxZADUUs7yxi
w0ggCfm/b8fmLFA4bxSQoKAzsTl0HWMk5IijFCfr1EG7EclhhgcsQUWCy4+nZfJi
g3JVTfI8cZhuvTeKfD3XSveOeBGDnf0TvK/zISaPMED8cfEHUhgB23EGdU9nnqtx
iv2KSHK+EO43MmrNXV1br+AwfVyunc0SI81MVPFZ2TeCvRcGwsnBjsU0SsXd4nVY
pPZ2EM/juqmAHsBkSWXI6H+hxL/SW3nK90qUY8ZNs09W0CkedEIyCFIE26BYVzD/
HjuAIUObo5DxCBei7hI9xF4ZzjU70/LRIszRJ3Khc2O5B2p+scx359Lrz4RH6djN
2+HOOfdvyxfVL/hU/EXOdgR8P0mccfSOe2R7o9BoeRUMEWxrhpE00o6KEn+AseCW
AqbVeidOUyHbpkVFTftLaRyXfAL8tZ/9ybSjyLAZRx1ryx56TkoYJ57bmJO4v4Ot
TZvsKYP2OQqmTHl5xHo3VwqyOXxQHL6ZVVE8EDm/QyqipsQUw9dFTs/yfPyq03PG
Qd4JcIRrFjOoNjrdCC5J4ZcRDHgzaZQ0dqXvG7Ru6EtLqS2AA9oyuoP0kkfKVOi6
u843KymFU9ktfUpu7TC+H+39bC2EGnR8rEwSFGZJVPipS98//dTQB2fkYBcsm1ug
JCoGUpcl7A76cKq852g9BvM29F+Y0X8H1hOWlWgMyDqFwYYB9gC8R7Zpld6dd99x
B1ZMYcOCq6swNvLcfJv86gedlN0tLt1h22d59XZID+XNvu8ECfkDC6XSUwDTKbN1
cg5DHBSr6ciQKEjhuYELdnWj52Y9jXWpFmMBtFPchxjooyjnCCL59Bu/FPqMnm71
OYVFEuQPNWSl1lG0MRYUtUVDbXPzNgZwFKrMFmOj7GAT54QqzfueKAXjFV3CFDHr
ktvcQj/Jj4Sw2k+3srCUvvTOFT+2hC9IrhILXTaiWuEFYx2+eYzp9zQqPMf8qJ7g
ay6f2IuqBljAe5/xYUp9NabT7oDyqJvCPaF+aMwt7+wzQjgD2pbkFAuTRtkyyZpf
VQhfWEcbjnfzN7+N2HAVUrHO+cdvAhd1zU/i74InFBp/5ZREmmFyoLN5K3MRMKZK
hKU15mAsc4ToVAbDRROP19FQWaaCj586Nx6WX52peVpM+h8Xt9e0690FaxKVU99A
kAqB9dPqsQSohrbDe+HroUwCqeg3AwJpjfg5SOtWgJaxXJULtfh7ilSjW7lsG80X
sIA1tzp8VDiim4EVnXHwhaCrdqoSkjVp19R62iA4yl88OYIU+9hBNfn/L5/YNZy2
uvv2a6zCSF86zbVFPr+khcSUIcD1afNs6/Zz8ZeTRAPUmN/chEweChhgCpyyjAbd
O7GhRORMCQ2o1mvRN3BMNYOJmdiHxP3Vb2Qxvtka9F4ZAqAa5V9d1MoCTqH2b2mR
18nWOq2KAPTA8w3Jl8mJDjXCAPrGRG1zeUjOyq59iBxArJ/pJm/bytqueeU1x+Vn
aFvaNFJb4bKzP/AHKzacNFy0KC0wuBfAZVKlfNyZdSFka5lhSo6VIRAqBFgpDebk
oPJ7o4XXN7wJ3lbfTxguVXPZN0tjH4Oj3gFpOJeRsv1eNpxerMfN1FbJBrmh1GY2
XJ/dNuC0XPgH0fZQWpcH3cD5vj9BFZAMR4EZ4MTw+PeYeFsVCl6f9MMC89ncxqt4
/JwVpB1boqa/WMDM06MsdTIucylXwoiBrQ0qXGR0KSjB8zkKO9m/YfPdrHGmxLDq
4dI4w7LHmMgYD1jfPxcFaSvI7Fl++2v0L9543KXVoDoXh3Fot1pYsCJGFTTUl2yj
S4l4UZ/buXwy/MH4DO6hyMrhOJDEH6UpeyMZtdvQZN4g+MXD5ZXq9wnrrqFIftsP
ap9zRfc6vXy7W4zmuF+mEGqbNmCh5PRWEkyR+7nHsyDCHNWinES6oPSph536zA0p
DdwFyZoJ/zXsIYIQJ7Hzzpt6k/IDz6JyDo1bZ2fhiNqV1DQuXWIrbqQwcSl+Na9q
DJLk58xOQf34S08GQaamOoFpjG8piiZDjRu4BBcICm/vceLCmihCaEBw5IiOf29i
NKfyAAwq8VRv3IS4cL8h+K7sX/3x8UQv0/h33iJBr7x9dR478iCgAgFxUOLqRzmU
1td/PqQPfhmPKAy2XTPmczjZyMAbJ2tlXMmYuG8gQXGM7RlimjE/2V3spFGIWm9F
8/kPiRLFriQxwAIS/psv0qCcdvltKhn/a0rD/n2iLzJpRuUAviW4d55GsAJOo0I2
5xC45C1ih1RYNl2fEElhBu8QCqo2hEMMG+ZvmMpRpQcqL+OpLtjRA+4FHAj4Fnqb
ktYiqyETmQVLu/2c8kQknLiIv0AEs3zA4+mwrnUEf0iG+rNM0g1Pm6WtWTcd6Tas
3L+6bIvkoFT9XcrivFmNbyDde1hakLwhTOpxNKlvNhO2cNFGs8MBOPHRmtR5wFVU
e3dSZDhMjMqfRmYEPqdmHHmQvRrYq25Tw7JnraACTC/cgdV0WUfpFn4Y/T74h6ny
PE1nV7+K7XZJfTmgFL2IslHppDqd92HDRWzfFgALqaUouUrVwFbnzV5NEGGhRJ0j
IkEqLhUabDI1K7bAU6mI7KWz/ichQRJne4CJLeuz1fZ2yIc9W+AupH+HY1ZLWXxz
N1RXuOHPFv/aF8FxApyqn9FnOx4hLkPti6PJbr68bbvntF+hWxJrChewncMV/Vfm
CudC0FtvqIQ7fxD2Hy67LY4YgbYuhZWpLN+rZOGU8xFirxvrHsiAmQ41qqNgqsrJ
jZbHn3xoCE1g6Q4vkktYSF+wNGsIDiAGVB0bCWf5VakywSMpTl38qsYEXQu3OJ7A
S8CtlBCwhPw2f4CZ7St6b8nXNIHgXRmyJ4cmDVnkUn+nih+7sHyR0xXMOLW/0TWS
ebcHizWr2u4B36Y8U/1Zxmntufmfur0vE84SkK4wukikj/MN7a2WLFrJm3Vc/Tib
jFE3V6EdW4wypXMLQ/p4cvJcNLRvH6+2OkwJ/b3jP8xj+7ADNumLs96SKefGKAN1
uX1Rrgs7N9ZAt7HAav0zG3zs+FxR7h0b3Hq31CcDIQs20pK4BCMZHcwLduRu5/vw
eEC5JjN+vqFIyX3PiCw1VdA92ZT/C4m5RYzpj4dnIkZYo9x0DSXGNh1VtH0yezC8
OOAcdPiMwJgy9aUC4NgLK3P9y6CwCAASrRdKStCXd2PxwQgUoqeYLfjI3JSqEjp0
aWzaN6Z0El+Am7i/ENUimnWcJZlyf0+8eCQQwvFV5mU3FmNK22cDIUoQc9iYq7ac
kvzQQlSR1NI9U5lEoR9gVkBix+ASgajCfp1xR8krIDTUheIuL4FAaVBNcTXEJYvg
jB9AM3zfxszp9UZ4ZPDGHqPvQawswkKFllnrAJoslv9BPJkYyJTA5Y6gU7TP6NdW
xs6x3jLvb5SP48pOjKmdrbsjWTt2FHMIiMoKC83tB5Z4B2X53OIDtXiisfVLaYYV
NM5TNl8p1d9ySdtGIQV90FMhk7q5VrGLYZchumrZXkOzHkTzYWZtFJisi0zrQob2
lco1JifoJHE7m3rMVsvRedw727fdE60/WV0XsNQLWZOuB5IG61keLJaNJbqy32SO
X+Cs/dihcfHuT8OFvSxVam2ayhKp+vU73trtZLCKS3JQuY2D0WG2aCgbCdNuHdxV
Lqn6qBstWukPU15UnGv8o5hJVG10gtRfjb3qUNF+WV8MK/urADbVr+31+pWgGzz3
BH+kgEmhJMbbclxJXXcDTdfn1H+x9yKet0Bs+8pq+OO+ctu1TOulvq6qUYOSHegy
tPTd1rG+8K2ZWos66fZLn1qVi0YKC79KSf6Y+iwSzGJzoUSG0Z2/me8OTA95gftG
BaBUdZfT0gLmmY8FqnSrAQAA/dQSt99/3YfHygmkX0NJh2j4XzwXdUE7m9/XCJl7
R8+u9cqcXFsV14GP/VQNb+8kg0IAi7WvCh6qpwEJKn5bsBpDIwSS2Co7A+zkqZh8
mUmsvBy42p17VOIZkjD6QR+Gx91am2us2Egk0bkp2Q8XTaZnwk+ps5zIyj+m9+0c
FxHu6/e3k/ZSlbom0tfDpe4Z5/B8zv/2nFIQcsO8eiZ4kNqfTMtudzFrjbF0uMjS
aWXVLJ8pfvqr+SxdioYQbReh2iIa5lk3YpznQuztcsgQJC/j0oUlCXJ8C4WM1yL/
4AmSVaGnWJGgrMsL4HoWHE0cFAGTiK8NjrPJ2Bjpdxwg0KBOOWU9C2/Vn2jhN5BO
k6B9fWxGeGkwnT+hERYQQYS0WVl3Y3nrfvaZk7zNSWkbfeVZZCD0ON2VClQCV5w1
iherzgbv4TQwccF+qO2hSGXwsMEJFN9K5/eVyBo0zgRt9/8qdY9JuOVSdbJE0p/C
hyqP+M4TweAfSudJTdBgdLRQjBmDrHh3hjNhCGvRFfIOaZIywyASgf7okOW1oEJj
T5SGbVlFAMnby94Lb+TgD69Q6doI8mwFg9CQvlQ5MBrRYlQZal014BtkeN3BDjOv
ej1/i/lsM7TrPPl1xD4+7lsjQk0K3ce59ZK2Aze4MtMmS3mnxCSQxOpAtsAuJ5L6
vohQiiIivCP1lcn7j88Yjss+I1/VETaTLrengSHG3NHtFS/NDeVfTjBIFFnjJ9eF
V1bh78tuOh4eHCTCkQxn+Bn87CvsMYvaI+/K9+lqJzkCNBtI7gKAtq00+7ThNAQo
t7WDTz2P8vun5AQjH1uD7hxNgBCJDs8TL2LaKmZFLB48kyHpwzZIIrYlrwQSA2JT
OFwwju4IhwfoGrTVQHQ9cdDQwnOfIcBo46CuIBMHgH7yRsWYMgKVoIK60yu1+QBH
tyjrmPglIEkQaT0LJB7vJBNFVtRjvK3uGPDGzars7Y3jiyqjkfVzz02rxNviBC8g
elExk+GK/5PgKkatsA2b2J9h59VMrBXp6kgiwinL17VxtvKuESOpoKzwYFlJ3H7b
3/Rzafxiiooq3hWtd5WMJkholamHrAHcj5CIUh7Wg/QVSeNCxcmpR6D/jWPiS63j
WX56pLY56LWQsozS8Zi7GZhxR4kNmGD/uFvsXbBnbCjfWhhOiWFgIEYIPb/gqjKr
TlghN5niNwmxt1TucrIRsbRZD9Y7fz9pqNBbPGijJTBytqqgGYoLdluDn+qqEiby
HFc2GdbJAjEKHzuAiNqzb3KXZu191pGZMxMuxjvFZ/a91fR5vEnvcZFG/ln7h5B9
gUSGWpBPqqMjaUG91GzH+ZU31wuQOos3+dJVxA0GUnRPKUtg3IPNhfVtk5qP+e+h
U/PiD4JrBShU+9FlZYbQ9Rw2SjCKoplM09mDoxyGitTLoc+dXLtWfjk0zoHK2Xu8
pajiWnWa8kXl+8R94BGQ6CvDeAB0OuY23m6/6BQuSwzugmutmF5Fo7i4ArDw1YFu
OhALC2HSNlCbCcUgsCtUTfnGoqznPeXzA/teN9Yj1TlWGc6W6E9hC4y9HKCAazLJ
W+A+4kes6cfP2FBuatP8VrAnrKLuL3A5LMIHZLsMDxgPx2688BSE0OH2+mrbYqBW
jVA0Uy4abbPXxVbjU6pJFiabVviWR+OYDvxYUbKe9rN/AaunIbBalsG6tEtgLSOr
ZcXYbkLM2nXU1wlOsY4LqSHgg5l+p1C1s4SAYoQMJz5QMDS+Wtr3FpdqeGYE8zPb
v2pxPnZVkSNLHlEILUsnGsewkN8lrX+StdolKmN+9Ul6R3kZ3UWFt8bKNTZRkvYp
q6ndxuFLhPre++Mn4UXxTX66f2bMFvguygIcaRBvvoofNnnLyT9RWeO+nsxkYtyG
oLi8BSfDvHKHKpPnBltbeJkqZQ4AmbFR7pYmmZO6zyJudGwOoxRUa3BMJhPgS/9N
v8795X+LX9/jQblB8lY9pDS0+nknhL3Nw8t04dVbQm/hdu78hJUKhGeIyCZlm9sM
uYZ6DzRGDHd4IyJa6ZNA2rr1E4861ekJJmD5JUcAsZ21s2S+lI9jT7GR7fCjjidx
jvo0g+Hek3UczM9bnWjqvag92778O4HnbDq//EIu2kpyTDXgknsclWOXNkr2MlzI
oHtTxmXpfS6Ix7w+iED8Xp31HejsfRql424DqZfosVGsR0qRQx1PvHTDWP8ebWoh
rUiTtolqiiMAqECCv1HcltTLSUv8OAwqWOHZEcK/2skHYTuxQMv//xijY2jpec2L
oZLPIR0EYY6B35smtreotTxUqpHekGK7dA7sSvNAO6R36gbOTO2X24T+PqzMxjZn
+qkUR8LpX4kDcR5gIAUzqHXAyCruKGEmGekIp3eE+GgOLgRIXKePtI08FsW3DJUV
H124v3Y7bWv6lzkG/5F3VGrBvcdG6/1NmVsRnH5bnHpGBBCKafaqnnxhBSA4JoS1
u6/W2RDjOk+xcjkOWb2AW/0MZx87fyr1uXuHMRPbWxvuV/xg/MwtbmTpQIJGA9Ye
L6Chronp6HOEXWx3Ww18U4J5y3olqXVKPzN5Fe4F8Sknbzhkh4nJ+0ledRAhmjSu
8O+R0pphBD7Iou82wQUrDjVz3Y6DQh6rd6tq/ZDObSH7t3kkGltU/gAAs1KT0BUh
9HeLe2f8PteLs2qvl/b6DfO3RfuqkmI/WJ4Ka2u8xqdcCDLjV8nLMxAc90D+n3Qd
h/QIGC+n58I4VBdrDjznx5cBqUddpHGH4sQq0+BohJrr2Cf4a5LIWJYuPGUfSvOy
EV15w0iM3oRPg3KB9/Va37TR5Za3GCgaOG+zVs7D6gwNr5H3p1wlHy6nlxDixmV5
PZh8flmVbcR/PO4iWDjGg0Zx9xIlNtgQvytvgFNQZLZneIQJhX6Co/EioJ92rZG4
nkKdcF8ZauWfRnxBGmmliFvQbv9M6lY5RUZQw/upYQEbUf2pOVSX7OpZc0B8ZCPq
qR1uANY4FAIi0OO+fLr0jkNSMkqo9t2T9N4t5kkEPQNNclnd8jALpFDRjIKtXq04
qmdfDlf1tQxt23rO8CpGppVG1t2dGJM9ruqOcvDyCGlZtGpK1AyaSq3JYePR0Yi1
M5ZIY9rjDy0m6MeHycRJ74R7INw5q4GPGCouCzWRZusLeUjwe6NOdo2ej7YI2BcG
7iEayf1+NV67yrHQsLyLwv7v+SX6bKnRNSfE6skNkOlfWw6chlzCevvRg931cVKA
EcaDJXO8RDwlTW7qpfp58o6lHgzxOtX5bdpU9zc6jkdJv8gFcELWEeflXmr4tHXd
OUJ5sS2dZqsNA05zzlUpJizEN6d3IUWW7xifVizoFAUqKKgbGYeQkRX6Ny8HD2GM
i/RbJXgrvJUDoxIYk2wyhUq+8fZv/WXk3dFyYWbPo9fp16e9SgNndgoxILXsS6al
b4qIk7RZOhJH04mxdVZ0OeT1TR4To+MswOxvBjcVWINOAIMZbfL+wGVIhdYyN4XU
DKNFkrYVGZDhrCerTPRTGcVp3ikheCOhCCfJtaSHCAr2G/o0cEtEiNYKtGwdMTJE
VQbHj1hmuDsT51SvqNh1yY7x6jJiAU8Ths/DDmH8DfAtnV/+S1Qef3v+TrjRNq6X
oocQ8Gi9tO8Niuvr83D6ohRNA8sSiYirvljvSpHyjFE13/eWNUdYBVteL7xXg8kl
cXVVqAEjKYKTrY29NZ/jts02aMnAke53aLmHIYiTZ5Ocp2UTUi2CT2jXdnlxXbSi
XvyyJGnR50UgnrhbKAREDPGZ0GreUTxfxAiJjbwwnLImgi6UbA8qs4NLX5cEoVjp
1AIaiObA9w1C0Vd99n3udYJ/zbIWqKMfHn5BCzbWVyHmipaXRziEMwwvDPsy4a8w
9IeZj/UrysF/eqpeS5UT/QJkRPV+/hLiPJP0nMwZsNOhq9DEmGLukoWuMJLyA/ph
Rc8mZu5rEtW6I6IVvCehrHfUat8aSQuvmHJNkHmah9etB9OiYJR0flDD77PcVL6p
WUJeet+CHl8d1r81ypDLSdhjVX2FIZTe56LDJ4i8caiz8Nl1XjI/RHiQip3ZrB54
axxwbN5IAJox4uuykOOZ5cR1PjHhBoFhDFIfOfnqz7rtcRZpIgivZgMfCqJ08NgY
BXsWg/KR4TmBeznGoG2dUWUxDxCJHpPXF7ARKKBJLwG3WJIXNibNb7o/fkqZE60i
sUhL13JURFpQcZU5fBHg97IXDgEjJwBJC4GWhGa4cc+OHBUj3p5sxOZ1iUp3CBHx
LkKbmCOCRsq6suCBHbLgIbQYJFGYsPpNMYp16v906yEvzwnVPUq+a2WdGNV2oj5j
F9GQ5Z7o3OtIpCOLOYVm+1+hJYEHZt3deY6xX9d8P1bnQ/KYcSYFuTTAlYlLvNP4
q6gjE7sikY1Mfzbfl/qbDza80YLyNTcrekWlnSjPCppDDsZwxpzVISC3tS+2rAxh
gHG6y+gkLDMHce1tya5yUewmt4stM1s7J20OCyQ/InyfTkT5WgPmB7NgI8ue8pUo
qr2P6dubd+rKWDbsTgfNECfthsOdwz7Bi10gFUtMHZ/TdKj3nFJouaojNQgY7k6K
tXreLdjH9fqa/6MOJaNne94Jn2SE/L4NijDas8QvRfWiL7We6E5bkW2ZUARFWAKm
p+sJt/LjumUDT5H44N4BJOliz4qGBMhTNB5yEhwfRwWokwHL15o65Ltb9RRXUYZn
v8I0vNaEf2Tx6C0f0QT79f56DbHzg0aLMjE42Ta1ICkgqRHy/J/69fVacxOPsjtw
Czk27FZ4i7+2O+/V3tYuk7unpR220WSYmlTd63oUANgFMZKiVLj9F24hYmfY5hPo
cP+xnmLlFLEtg8bN3qxIs0nfR9nmCg0NdtNncH4R8DC7d35r2aXVer+HvfVeHPUA
1N0LNM0eWWeXBoyxDhZP16QXLU4hz34PX9XI+ArKUkXP503J2dIRN8Cbvwo1c/7a
znatO5XTGquSjCrgAn1B9fRF++88pc6qbnPP26+pGGhEspsTP9404C4qqzKyeHyG
Wtz0Oycowc5DpGl38aQcS59C1il+gctBo7DZt6FF3VqTum1LYO2o5ELYdqnLasz9
lScLz1k3a/d3hoiUN/xFpbVJIJvcBKhNJhUJlG3B4fke7VQb2QnJFu0cAXHKHp09
3Mh5vfKIlnqbnDsP5kfQ3lKoNhEFJBGUTICNgR0OXsVWBuhrxJTFFG0JnOZ8HLeA
LwvaRntGkfHYKDMqhWweYPb4fuDUoGTatsnvw4E2WbLTN2fS35ktigSckyPTNjTb
tCRptQLjEu9zmVNAJRdd5vAmEfYjKzox61U9diOYR7nu+Sm5ozxW1ils5c/mxrfS
mQWTwQRzXfGUWKuNm5sutSfIll+USt93ZCGlZqoyFruWmVm5JECi9qXh9x0eloXJ
OjCapP6vXN8cqZ9POMJbzAqu6Y9G+LjxrMNZBy223xGzW+Rvtwtp5Tr44JdqmnI+
cMk4M+53G/QYXVTs8pcivkxO9l33qALl9N6olSXkdPdYM13NWN84B4NapcU96nhT
aPyMCE03EfYRjfwXnaphSpZuVuPpXz8BT6XaoaazZtI8xoDa0ECJWY2JW6GsJzX5
cmmB4H3eYWXeMN2y5vPwAGPPkPZpTvKPi9EYRR7eh/D8Xq39d5NkYtyyBhHiQVka
jlF57bcBEK9IWM81K8MNB6lSpXcofcAqDu836UhpAV53+UbkQMNe89K+6axadWx/
B/R+eNmR9udz2gmfi80U401wx8f57utR8Dt0ZOuAQYeUWLKllsv0rIAP1qO0rsjP
qxo2wPK6wn/n+8ohcjAwMjfMCA31V/Cb2Lx3/W63D1md8kj9iWlzKfv8xWwtiqmF
o6eoxyXfzAwtIEs5Negj+TrB3su7FrCtpz8U/VBahV5gX2XaHvfni2WJX34XaweH
FOel6LJl+YNEpISV/ebgJnR1BcVDxHHDjh1DNpHMgp5+eHfRGItJkwc9ImJpoNMe
Nj6NIUeP61Mh8MyAvXJJm7shdh5NSRNIgX3oEI4Ni2bQDub6nqa4ZLzVQ0+CjiGN
a5VFBeqSwdzQaM1U/e9QPlxVmrvON2ndr4izJtUr5WJtaSCfrzXAZk6znRYXpA2F
3RMO25hGTTUQksLCRNr7Cbruooau+2E9oEPwGORH+5Jybg99hFWgAci5OBwHdF10
HH41Njg/qZEWd772xHNKwyfPkDhax6My1VL/wKHcLecXgh1DORyyHaSVY1e50b4I
ftGpQs7/3pA0siiEJNeTPMxMMKj33WSzWw7yZsaox7FZjULiL75UBX0OzK7pj3a/
Aqa9qhNwmLUjJb3WBhx6FYd5eju60opyuyZmis7o8I8EyjbA+DUKbMueF4fbalGy
YUs6VzWJMcSZY4cHstFFj7JugdszBA+eJKaLKpGDBGvicP5tcPEiPB413A4e4Yv4
h7qowaz0Qmb/Up/TDjTyeDY7HIB09xlnw51PxhX941SsBjDXnAh3h/Dxu6O0iDLB
lMA891wRs2vCIrQ0vOPrAhxJ1dP0pkSjacNZhCUMhy253o2wcHGoPrEdJSBCEKd4
N88K6uRs76iUNEtsRSYhn+rN52ZSCsfszwA/r4hkHJOIir9pdiXI/sEvxKzsUF2d
MpZX43smKvCQcFBktfsHSuN/00EWI1Gk2CUB3EZME3GKxaxycdCWLICfVOaqQBUx
ePyfZSAXV+uKpem/gcxLXTdPqmKg/+9mhPq6zTkVzZ7QcMdYfAxvnH2YlXyISMPW
SVo91KV2vrKuU1wthVsPOiOmUQtLJHL9mT7hJhDbH7LUAEw5xTxtPNn1tij6POo9
mxagHOrfekc+F7rRaK1fWXQHmA+JVRlb/Sktm+aOq5s8EEhVJNpVXp/ABiV4/znE
0kQcG3uq+nrmeE9W2nDyA4qHTNUSVjyruqRIptJTEM++ADtbTqiObItKb6vhvOEh
ZA1C70QdSXo3ZVlbSlU/YHfUvKLrEJpIG4EJgSeOySsdhNQRce3bZOKlmg3kIg6j
k9hBbAwz2qdnDaDARfOfPNODGC6tBk25ealE+HKkWUr6/kRBjR0XoERRYCXOmnvs
vP71vIcL/3B0YkonXKxtl2rnQWygACxwDdUJgcqQxHDTf1Vl7cIF2JWTJMPr8JkG
nxHmp/amUI1YKwL8EwnD/DvUn+dV1l8g/4WN/SMNU3kRp8MnRm3GauqQaa9crylv
xwA3eiu9fF+T1Y5GkTQf3bLw7RCTxMD7FIUL4mpkm3qsiw+4VuYgIOWXX50/fKvY
XY+SbGaaQpzcF4R9S+tAggju1uxgZiej4ZHbTlMqLXH7e5N5787zRjdndjD1bYeQ
JxVdkuzHcnr3x6i4z5O7HbDkqsR3dhadOBZYQAn/J1bBIXmtPtvyX2VyquAtIWVj
mDYBGba3r5vKXgeSF1+J5Qro4L7zPTKepqlMfjgDewupMSS/3ZBM6QAzrqKnCyv9
p3y4gAM0zqJj+TGw2703MhnS8d7Mg2CZ9SNyA5+pVCh2jVKk1FaxSHN6Eul0SGtO
1gr16gZqIYspvDMyEjjOxkDqNh6UKBYvSUWtdHx/AR+fKzDSLjOIjRNGGuzQD6bo
mMHlbLSALzJlspbwkpoCKWBiGeSb0uaLogFxQCzD+qqwqnaEq+fuyJKPA9EDbNBF
Du8t2oIQjwiscMW6zGQZ4tOwQoQwD+z6V7vijB//+Z+YSVUaSqTL7e1CY6ixSbYj
kg83kTnpR+OMyqlqATLD8yH+omHzusu+2Yb220e6aWq7u081x+mhZh37FDzVg5SQ
MUPu+aIMgg3VYLF6zS5a85TYMeEvws1SV3iVFkRC3QhJJ0AfUQF/yX7BG3ZtsA2D
wJEty8Dh6NHsRnm1p9xwfy/SpDNh7HcV1AeEj4Dg7h+rdxfuYpdKhhfsctk6q70f
UzUYrcwb96UKEy2qOdQd1QD/wlyiJmDoxOXRi/Fq7Q1BGmE84cmpUrwVwopn7vJQ
j+8VuBWp09ci0UK7nAryuMMCOLza9MsEERtTltx4MN/LEcd6J+OAvNHCBRSDZolz
HWfg+Cqkbfs112q2uRwjJ73CSvmg0QyH9bEqTNpMLRHAejyLKPxrvO9TsH0RaU4B
CAQ0fgO8rkpLm8+yYdld9kjmmhSo0X+TX6xwW9C3LAZ3pyO4EJKBajMCwneV7dhU
nYiS/oVD3HEifqkUWg+xKiXFF02y9KGWWD2oOQCsv588mly6DmY4VDIr75mxgW57
/ZfIs0lrTXzsYJlOY6LdW90xuB77RmCKb3dJjym/lWbfxFWvDlxlCIXGDkHijddm
qdE8FHI+f5/xTe5lhT6XeEJzDhR0znHvSv/Flu8hOjIR92MwwbeKE4zfXgZynxsh
avbT/BUGJmSyboG2IOx/negXQjF6gOzUwoap8XOgLp+UUjva5wkz3ZPPBgwD76Qs
jNH8hLNF+oC5x16XaKEWzfxxrK79SNpI2buB+bKsjgcOiCo1cLzEGJefGZtGCFeT
SPMtX4FpYFbOQp+IMaJ8HW5EY9n9xa6R/cUvFqmEiZxcs4PRjJc02Dt1N/UvrPXf
g2BoFyJ8Y2mAkFbSe/TyMuxI3HjyUwHMwHmGKedl8NydoMflfkUZz5XHrRcIt7p+
lxNmal5PYGPEx+ifiChW24ZN0uzBj6NVCrabZBvU7r6jSPWSs7dHBJjSdTNPYFHe
jMXcT+Mlud4A01brgZVWLMNDadfROYcfGCc/PyYBLq32yPYfBbHDJLX3yRCExghs
wpaKVkjTbbk66iKCyUA1PNkPrCvMhEsrotqCxvKqnwB7qDOdLX7dNL14R4zFLXlJ
LxH7XC+6xnw6LXSQG3hcjCJPRM8YUbL6Wns6VekDVJa+2NOzP4NvRTtsFG/cjCcv
CezgW3qAzGasA8eqniV9LeRzGhk+F7vUS5B0MqYUzxeuGJ6kXU/LFfKivy6TK0tI
eL1r4ACod26TOUmk05XS1FzFUKUrIsvbc1xUHRCeCZ8vCbGB5tGhpW/mEPPfjiqg
WJqlmuzXNh55XVbGS2mmVbcyerImJFI58km4F9j2pYgMEfGN1VHSOwT/2TGqWVJL
mQ9yYNUp1cE9MyZHUQMlEVbmh+2+Lvfxao6Axvq1Bp+lPgGDSE/KISTsT7uxCp06
6sOrObY5cb5rz1OBsLklqq8Vy8KlPSZzaOb2WRZPHQjWIcJg6mMMpq+pKBVuGL3g
lBdsH8WClgxUIgL0MtFQTYcXHrZbnbnUHJDcIeymFUMgKq2nHEVPdvV8pKH9RB3h
kVGWQd5gztPp782oG2psFxOLa53tTXdQ9z8v5YMZMMCthpON7igDDGVp7c4u/iIu
EizlYPXSEd5uIcJyO1fCB7rxwEtvVq5gvB5OVpVNNC6EVBKzhOhYT6Ob4AUJ3dHp
rT5lpqe2zFURAdXue6GxNyJWuYOrDlomyWdyEznydgWPEcWDMY1aQORJHnH5i7bP
6GfR3Y638nYqHSSIDR49aoWfV/4+YEuPVd+pOJmqkCPvB9zFikABn/je/lkx3881
SRbUKhT2KoXhX+wE2y4jJZ+beQEIiFIx+T3N0vCAakEt25ASfn7+TYGCK9IfAL7L
XyUXdPYu3rohEGGXoRr/xI6ko4hVjAGWm0JH9BSGaB7v9Xo2h+WNNXpbCOoFo6tM
wrqLlIbDmlxSXzgNpPZSzf2NMAFgBbcZdu/mMXQQPBZis3hUQHYy62spMS3SERhf
iQpT5H8/Jeo/ZkulNFnDfhP5M3cjuBF8U3GkaIIqnfj2TLm1M5l5NLOxpWwNSGPS
GH+5MBGURYASzVyiw3kKttYdXEdc6SL8/0t7XK6BbeqP+Ex0T40qPNU2copdif2j
08HktCU+B9lhKILDuTsWCHkDkB8J3m9XPXdMB0smiAzQZ1xPcz4EGjTgiYzL/FIY
VMrTufx9GxEii9/YbIZyDTouz4npVzkQS6xQvBukBeC8BtBigFDPQ4BU3A7BvHI0
S1wMKpFzTTqzJHbvgkRiLsv2oU2Kdhrc3Znkw4qKqaP6GcxJ6+hVSfuDVTWzg8AP
aguWIpjsRGcGDOTPDE7m1rtD7hDV49cYkHzltTfNvNFQVXkeaXZ8K73SJM+2yCuh
L9PzG9RgMtsjtpTGyFYPICM8QNLAG/DoQW+ZH0hkIJfYIn15mtBvSzpRqgKJDs1q
XBiJfsxJRoVPsVbGs1b2336t84hwD3U2Qs5KPGP/fPZMT7s3JZV5nbs8rfnTpZKx
YRnYt+fIUplvsVWNTRJ//6/JN2dBEVlOOn3x7bMnhQq/XtXOCnCNbEWc4aOGxH/D
6BOZu3xWJ31Ci4xq2QMCPHnrPb77+X10mRFRziRdBZ6xotryaIwHTWUGWfrqNwDO
DNDKUWXTMUS+ccj1KoiFxKMBRgrgKt+hDTfEcEXE9UgsfTrc39NecVSb03v03VQn
zM4ZpQFctgjI2PTjyNVzGbxWufphl5W7pZHkDjaZZ1M1H5EWz9npAESU2MaBJFyR
zbq15kwFy3AVshl/0+494IGtWJuSe6KBtFuTkeSfr0VBNY3Dj//IGeOhsHRPL0xT
zBSf4orkYpjBuQm0mefOts01aBB0qbZ6i1ai0fAb8WWvsE49Hf/LR7CyndG7jRs9
T6plw5MMSwIPs+6s/faubCsm87ViyvI8ueuy9YKO70JZOwlfS03xwiDN5tTfQNXr
km0SPOViz3d8awdimyTU6zRly81MGCmkZ4aG0I63Pb0bqrQWIrLcgJY6WzxWl217
6dmNle/9SG6+CqKrNx53k7YzrPZ8HuOzIGfYGBKzQJtpXJDzF531z3jQ8eWt9m/P
iFs66YZqCWH9xuDzoI7IRgv1cjf301M7wYtl9qLIRV5en6DhBbACRm7AhnzSMPY3
h3qU0XX1oagtbvKUruaipy10gk2kLxF1T+f0bgFpsIMkkysYi+IFcSiXdUu2MRR5
2vVtuerNVLnpwGAZqfZQfZH/fUGu1KU5CJLgFtQBrMGrLbuEYYcifDSw4lzkHjgV
zwSQrJ0tLMoIDrrN1sI95Ik/bBbZMLJTx5tACuAkL5gEI+uQUyGZGb1aEnVN/GFD
XPu9Hv4nbQVYCNaSt+xSawHgdak0GX1t8O9rEWE3SEufvRNk21G7YRK1hdXU89of
7xBod3vs3g+1vwkvQ5Cjli4mT0kPCe6IDuWX5rQ6vISub8FpSfRGNFRUY12ozYx9
9QdSJLoMrjRAOTLtPI1jBiECpkm2yTDzhNw6orta7RtNUuMThw5wOK+aFAreUknk
CJ+ydKleuTiLZTZv4LCmPtoUlFJrdwJHs8yFpnwo6T/SEHsx+l9DyKV0ZSbYw+aM
VmHr2igh0M2Z56GrxW62X27SuNKIp8IM8+aUm731s4xZmWE24ysVG38vepU7AxbZ
6qjPIefPDxfv36tUEK62xMlHnel1plS1O6a8iD075daY7Ej5gkkGw5AckHPSR869
XGixfDGTZteeN/wHAgZmNgkFISobiJ86qtxIn5bnJ6z1cy9xWvOEQMH+/tHg4rYS
MJWjcmBCiTtS99e1gN0hXCxCcJOdQCsj584MAY+F+edInk9iHrXorGhsJ+9tB4d2
O49aps9WNCRETkm5M4hwfpa4oSrJN58bPVjTHvXmKfeMyMuVWGa+p15J4Y7Ij/mU
TXpSEBuj6Swyc6b3VR37rc1Iau1cC74YZO6D6LrWYGR3CuxA7Wha9aswd3NjFCzb
Hk/bYm7akd9Hq81u3n8qKuzyrEtciBk0YQsIKnDhQk3UFW56QcQ8t4RpOpZWc6Mz
itUNM7RXbLFkgg8a0EVW6VTOCMdG5ZhPz+T2OGOOvOHLKWWLHNuekXeDP4csz1rh
M8i87rOf9WUppD/yNXQqMd61ZrfmB/GEDQvweiW/LZQZFuhDVsLp146oa6HgAkFx
jUsClfraVfPnhhRORbtcCRwGHH7PimDIk/Rkani7SdrScCF7VfSxZxKOlmcjnTsP
KddXXjERDseondWtMYpAjx1J986be8sU6aAU5RNKpQmaG+aEMz+kmGeh5PQ0QVgD
9NE4np2fWyfbDlJmQBjTvnNWw+kjPj/LpDorT+MdhV3GK+S8o3NyMjcTlNV9njCt
Fy7RX2Rku3828aNncLIP8Zn4010QReZHwIfUrDTBqkKRIlmhYbrAleF+hF8NbuYf
rfA4LNQeqVq3YijOhsFpESEJsteDJjTRB4eq4uUt3iKGj6JQhcdMPyMR0ya0UBEf
3IaqpOvnZaor6uZ0RWOvR5rdZOoqp2SpeygWxtNa1eppDES1i43A71+l9+HtwiW4
SLRraqKMmMj2pEupZyrxFIpl1pZCmlhl/mQwfIHvim10nro/H+2zEwjioxDTm/81
IRX3Moe5DwbPD8eDJcwgT2vsJ1+CbH3bxQVUEhK2OkrfEc3vXBJ+RFkWWeKprp5O
KH0Ji16XYweO/xnO28FpBOeFfyyAwHEvd5nV2MordXzY747ztE/vH6BOsDY+4CQ2
IliTMFJzkwUeVLvhPFTA8dxP1xAW1wIm+mIpk4wZPa86pmL7bUodIqSj8NiZwgew
KufXstJTAVav4R/RfScPy66GYyMA+QqHGJpgCzWceMCM2xXkM0ogrXouUO18lLnK
bWEqETT1hikn5iq7To/7fFrGAwPLEhEWG5DSOMZKiKPu9J2UmvZabDMAvHl4GPnM
ucPQtn68ZfKRzPT7Xz/KdvP1MpW7GLIoju06JJbqPaqy2QS8diN/NrbDdIwMOLhY
UT+HsGQ4TECo/1NjpXuJOtiv4aiSAZP9QEzoNrTcAhUi5UjVOcssQiwTFeYUujp9
UxmcBuQIJ4YqGZAYfJqqBVdVBGFKOv0PeYc6xyrs3ErKrJV7SUJymziCo60GR0L5
kKZc4YYwIXLrHOEmwvCkIpH9jwLZDppDzjzK/r5Cnhq28Q9SdUgiV3yQySWy+Rlj
UpXkTWA50y8+3rQr9gG9iUiVEs2lvApVZ62y2DIEahmCgCWlerxurWQ45aAlTTiJ
FLRhRn2Zf9d3u0tkg4ZP1QiQ64B8g7YoosqNvsjvAKipA67PX2H9Im15IFcIuZVD
G8P2MFTrM0wAQFN44H0jhXPFA3IpzhwoZWZ3O6hd+AmXUQke4/TniYbmwE8SwiCv
ssY+Xa4A5o9YMXNTe20SGFoZT4xKInvRKE6BSlWpoJC6KsPDiLwAvdy0gnsG3QKP
t2fh1j3y+zZ4cO0JUXbKBR2ju7dxF3Qo5sYNNTgy7JfEP4mmwr9EwU7d5plCIB4k
BQLW+qW5sk1sLtiF9nm5d4cOmiiyeR4kEUd+n4XgDyzjb0tI6yvc16TXMswUiu96
QiZG9JsKA9T6ZbyZJX5LgTJToBQL8A4UQiQOTiF3t/XwCLttvjSfXSW3+wJsZl4O
lpeimZHflK7qysyKFcCJd36syDfOW/gfE5S70GK/G2c5Tq8vXkZC+nXzPwIaBqhS
5do4EoWYFz+FAbuuA2UkC7FKvIxM4g2XAR+wEgecxodCUDq0kmxGePeeFpaJKOTm
wqA0WCrSpapzxu4o8Jn+uGEz0Qz4g6Phw014nclU+CwWMVpqokDPXP2+0FcMC6SA
16lt5Evfi9W1LaUHVnAc7qIRPItRl3N0luFyDXGSDmQAPwxKgy3UswnP0QPfnAt/
63rEtf2PETSZZblAwAv7XIuq+udBk7kQJ3oL4TvDdx11NVH5KwAXOIsniJ1lZFOd
W0ZDHlRPkfA1S6vU3psiHQPQqEa07CXkns8LL/UN3FuvIgDsSlKsipy0mp0ecxXM
CAAHPj5moduNCwPE8sFqkOoFeTWGBJkw4YXRuDoB3mEps583QxTqvG3yaUmtmOnI
8nO35xFEEp0ZEtQFsdsHYUKCLFD5R13YADWDtMhylE8Fxd7upuYL2fzFMTAl4T9I
ygPckRGeIkasibPOzFC4fISUGQSTasw66wBIgUeODZBl5MDo9sYlixfdDTYedn0I
GfJEeiHIYwVlEhl0qvyOv0hySrpfdqDHEF40raLEOulpkmzOUH6T61ZEerBu1www
A4qG8pHEim4bkbf5SJNwXmv/SDsoFcqb7XQVhWSQK4y7X3F8cBFNbSMT7phDMcT/
XGSMaGeILZrrobXh1Bodlrk3shCifPBgFwv8NRSPeKr1dLGvxg96Uy97Q8oVplvJ
951Sw4hbxC9t9OuIAB6lmR0cxEw/CMuPEmWaLux4mrIuqJssh2w2dmxrYPrJNT64
DDsxIOohrkC1bw+/5hZkOSrYGQdysI2sl141dDofj0ixZinExRZnnQYn/Ml/B2u2
b1vSdQalkudDNEhCB5KqbYIljHMMzI6LNiYbAldeeJz6Sbh28mt4QQDaylJ7m6zJ
W2rGKMx6R1vstoY/WV72C/Ko/FZLyBpE8JWk0w4lI0/OwLswDAVOTEdMEhzhSlfb
W98UZ+CE90F174SxdtQ/d/CpAr694XP90KPA1WH3fEOVV+jxkYH99lor8sqFP/wv
oWQz2XMOj8bOVlwV1U54wUSDuabmNkD3qnbmUsLRNbixN5KmvwH0vdWUvxR4QzQ0
D4RdmemPt9nGjIntQ9lC2Wwurh2p0gO3HjVKjf4ILmGa5EwaW2k+cUswYWqF7Ci7
37ElSaDjDSBB71GYkPhB22ZaTuwxV93nmeX5V8AO2aVZZ7lPUerfCekU7h/oMSq1
TQ60eUqgWW1JRXDaIDLthu/XssNfafK0xta1j6UyMMDVLBiA2OW8rJ+hseQGOJMx
ENBi4J8Sv2BA+Bn2AFveuZ7fV+hAt/nDWOv/WUa8ZeX6P9ZgmuKVqdRqlqkw/rMM
xRSJR59jyWnR9TTG3dAEqvfVqcsmVDUzoktLYsf/R01+G9V3DJJqdKEIIpuhR6dZ
tvQqpumLmTc9Fq1IuZVpWZHHBdjRPCFBlWa653vzL8Y+/d8LU3pTzEaf8cEYwzas
293AdvKZEA4tk8cw6r6V+04EZENQvI3EA/+b51b2CXtJqmsJqIVNq+HEtwh41zpU
TMJnH7+ks6S3Pfqo+LLovGW+IF3DeMlpzybliR+kSSzkrZHpK26Quc3g7XBeAG2v
9tuer/HxsttclQiG73lmaYtKEhzqjrANm1pFnfm2KhrB9vqcDzCQETFRxal7FfF9
zaUu5epzbU7vgH5L0pVlpdVVo0QlCeP8hgfxqAYFCI5JO4XF0nBTGPBGoMGlVIkW
4M+2B0194jHtJr6RURKBEslTYREOov5qZqwo1EjuJH/TnFiXyVdaAFTmPD2UWWvD
OrLwWF4HTEWQYkcpxN2hM9V9Vqez/z8T9tvYLYRlOjR8Jq8EmZwpe3tEZfUJ15+n
ih3fgdmIWZ9C8OzpYsduVmfm8DC4rNvMi0hrJEytWg2a1wcyp72FzAYo4WlINn83
gRRQNP4jZG0s6OoNm3xqO6AVN9XVjAx1ldUU7666ZsBAcxriOQPXPfaC14bdk60O
rXeyRcoQIUibkruDFIay7KmFpIhmcKZGXAgg2yehB9p3LujLYUhHDL3TstPRNLhj
EqAJsfqwG0rufbFGuf/Q8KcQsqMCSCDn/D/oGHmQ3Lq4QmpmL55RrV9vM0kBgn7M
tgRLeac3NZqvPpG6QiMglT6szRV0NjL1+vMGkZws59NSzWWdQthBGgLqkaOenQYV
Ll6+WI6dNuCvHJGncn8jN8sD94tnO4HyogG2y8sgzTHM7T3ZE00i4MjOJxxNwTZM
9IviVljAQLwCB6Y5VCJtqxNv8FBaqczaCynVTQ9iQbSYFmneGvdxGNY1bhATm3ds
6N4plYdR31Dgk3zETIpWhZlj5ezs1ibNIw5JWtLwN5gDOinaamkNeKtTSygc66Qv
Ks18CLgC9j/3wf+KCoK+/dkJU3MwpMaNvB+3WKTGS1OuxJ1cQwrrlT6Y1hqoN5hJ
oQ3WyMQWW/oEWGfdt6OcFS/Ej7+SZ4n6r5ZP6xi4kIuOI9KAYRj0yjOlFIasLxDH
xpceIr3jzjxA6Idv+Yjl5NKK/JBgo9ASll2ICm/s5sZmJKdkVXO93u1sC1IOIoDY
TWMPoEB2oWIVDep0s4uHujo6VkF4zhtnrxscPM56nxgV1HUIGgOJowHHuk5lFlhM
SyZHciF+UkJFjJ1bJVHwk9ZbBZq0xecvzSrT0Aw93JUd7Y/znrXgnAZLAG+23nYD
CJifuBCP+OUnsxZw5XBnjqRFDpAp3ckNZxVpXhtZnHamEA30YHk9eR/MPX8CK8iN
+tYwXH4y+BFemELvxJcNk8U6I/07IxEWG1sbWc8EwHxEelW0XMJH3NTk4OlC9yYg
EXUzaEcSy04SV1Z850SKxaLwxKFOYYPbZCkhIt5MF765ToD9LPKywavwMgUxufCi
n+JX1eWeuVdlm1VZX7rfcYgjq2e1koYCslg9QS7M6WV/Oki4XIr+xHkPfalpova1
5SDacmP5mgpUkVkLLkMTwMW41m6gRYwALSNFVY5kruyUb+jS7It2Ug6Ra/Kw6Lh7
3jHZ2q9KP8E97MFkBh+7EMffAIe75VTMei431baFAShbDebatxgNS8c1NpKWSvrq
i8eX3bFa14XBbvhZ2mJ4KkYRQ/jKPUPWBPKsG29ICWUjs1dP0vOlVm4PB4Wgpjvx
G8qEFpv/MaWHx3DQEN4wIJZBIMUUKiB0k2A4+UBxGYK5AZN+Qlt/LYRnYTRsJZ2e
JqQsNX/itWxUxHocUaN+SeSszsRfCvrWhq5xLx2GBaRYBIE/q7MTJ+B7IrVRbZFr
7haMBaJf9afTlLeG659Md+/KTvU38//gdRVaPdEiOmfjAxDDxuMKKI2bLXlOaGiL
Df9HSvuCNzcxRu8P04I/QWRirarOiRz3WwIqEXYk94AKmVmF3yrKdvjXTLtG3rO3
mAJ83uBA/gwDTmIjl/8wDrN++pOmhsw7qrUlXUZOVPYlEGmfaS6CFc3b91HAcj3Q
5VvtsZOsGJ/4u8HVkiSHb7t9UyUwjtQifNjcppEHhuUHRta8Qmrmlme1gfWYL75L
DnwwQG2xXA+09DcDn48O2J2qVRrSnIQ01SevAuWPVfD9ujDBdVaGAsAurjmWM1GF
b18DQ4TGloWypq7kVKilj/PRd/WxMrrte84guHlOVNVcExaJRBxafj4Dd/ltPgi7
ZG5e+dzWiZ6qIQLzJt5mzV3ZwDkbIcg8LWIij9ajPoc7xWEWMsGhJCrjMbFEwVSS
6T67tEE4dzgjdi8tHjcIjJnAb4iBjf2sbBVHv+96eTcDjn4ztRTfNJYiKZNG2YsH
tqCT5p45To2zHYRzcU6+rdXpBCwvs+InbZXzUUVZf69VQFtjrUVV6nF8ZzKy/NuD
bhcsP62CEVsUO/0ci3BhJilLkc/CpxuH9XXuLdomNJqJaFUhK1dtA+LsCmnjj9cX
46pCtxzqP6KqZmp0DY41hOgD65BASTkFst1mvn6KAzDDn4tuF16B9s4lcjxpgxG6
qhcDH1Fn8jglxW4in8kOivBOakTq52SIApvGxNtJGiRJxOM3F/GUypXv/qgifBfy
FPV6UtX/c8GItEbNMLD0JeYVKJp3cgr4Ttzrmjc+GW3yUrkg22/x2V/4+3M/cvmX
tgd0XZBGVUnGiGOteZyXGPSNTUux15yM0vMnaZnKPyk/Uf+wGd4KAWxnobdy6/ZF
PCgvXHRCgs/9E8gRvdV9KTdjXzp01FCEz5mvYxA+KT3oQ0qH8DjP0kiOrM8CBdZo
nodHYeRBFG3LKPVV/MCx8HYt13HKcLhReogCi7WKAJNTJrEYyJgFiA4ZIIEmWiWa
D+apf9WNgTbf+sR41s/bNXQLnbS0d4CTS8Vw9A0A98skaqGtlaV2OA4xTVyIzdvL
utXDmSiH1vAzjvw2E10PJUs9Ykz4zlSB+Ef326NcV1Zs1UFo8j7DzfY029/bCBDC
bUSCmKHR8dfmqaQ4GfIkrW0FHK0+/yUJwMfPJCKevsERTHsuR7Lzq0NxOxeLFK7Y
1vk1QItrrjHocq05CMbNnZ3uMedhWZaqqmZrf2m2NKU2FMgjcCp6FW3Q4Jm6LgNo
loyUgzcAhQflIW+jIxJrSWL05SD///+zdLbhJMvZWeXsGNoxifr3tMuyY9+4opKh
82UkPbo3UiW2thIzfh4Du38VljSzO83qNpRhU1iSAGHWJxwzZtmXO1bK9pLKdWvL
JJ+jntTQWvPfzMVXV1Qt8UEGPD1sXRn+6jf8gmyify3xuLM/1KeU+3CcziWHa2ro
cien/DEbw6C2j8LqNRTEa0eKhSrZIu8MJQwqIWL2OnDrtP5R7uEkd8QpDzf9XsQE
zH1dxz/iBYlEli+Fi0nP8Yv73RS3jDw73HU4w66uqI+vdgE2Vu3w8CDAdAEsRoa0
x7BWKd7F0vso/ZkwpunE4oFXIT2pfv9/3jnc1F8PrU58+UwHv5uU45PFR9givmBj
r5Zg+5KKUY7EYdG60uyVcUZcFNGpg1BAt/yF3xr62ZbMfXBN97eRverrRjVbCs4F
GBobspf6jtuv/drUMxxqt7mxU2fa899C3S8sMc+b8M9YeQWmhqHcmxXMQ+tBJ02x
fImQTh5RK9s9ZD0e/8vMHbq/Cx9mxVdzlpnjTyK4VIPczxZaQdUQtIVuUPU45aTJ
qQ6Kl7wwAjBQ0pFvTCx98tdqLKEzKhrmlG8ui5C3vLmPma5slywQVwIQZoq2YwPx
tF25W3SrmkToKXahB+0b9FUS/+DGGwtawSEr52rYyeyw691UX9Ssb3I1hhZSsC4f
dvM4PDiOhkQvaRGe4ID2/d9IeiDK3MF0Ct5o8n4RlmoXonA+M/1/GUn8T314XABE
HtDU2DxKP+G32DywFStkwkZ9Zu2s20FEZIZu8la0jjNiqwU/Sl/pcznqLh6LCayc
O/eH37FmXhIO2AhKiaew5EEAtHTwK/yiEpq7a5zMJxYClgzkr3WP8rqZwTVSw5KK
6yW/BYDDCNFb/O99XctuhEvJO2T2oMQ1C+5ynXcekTvhBSuXCXHDYwPy03+eWvLZ
u1yHUPvLWWUbTUEdRAmGyBxntRCDTHNsAoT/5B5a20v7tND3gRu/9O2HZoKlfjWy
U001NRsuWO4ceuxHbSmk8yb9wHSYBL1ovWuE6hSeINrUr7WPx6EDBlP34x4IUcrN
SV7azsYOi6tis07+tYrLnxWXEzbW6ULU0g3W/2SChlzl1ICNvHT864p9RSCgAl/x
vR4UlIkD6vXQbBpgOv9Cm78CKSUz80CVC8SUI+Jesl+S/Z9XklR+zVnIIi83IB+M
TAr2l0uZeSZOnCxBrLdHHxY1HMuY45nKg4RQBo5SyQyCSH4BbApRyWRUYsde2Gx1
DMkM22Lz8zR39aGRBLIL54buSFhdWsYPTsGZ8OmS88x2hVXhP2T8Bagy1RrFiFvV
WxPuLjV2/LjQcgeqBIpIuKTbO4WDUQTGMEkkO5/CsvKw+3QhvHNOt+Zr/o1Df1jg
jbITjA2wE9EVCVl0xyiblj51nbhuq8Bgs4M/+bZ+T2C1VXcP2DnmYqtbijd8+5uB
smKboGJoekvrE3oILwcQGwvGYSRrvuqJC60+BFoMObM1XP7xHTgvdLtI56XHLZyw
AeCiZwfgvIUg+i1eLoNFChUA2Ye+NHSBvYedK1vLfR1p8QRUWQw7D0BRo6o2x4BJ
QpxYUB256Qw3YWKGb+r7JuI5RjqMr6BVo/dDl6inAND32al0cFtMCIyfAPcZlFdu
ieoIDNzRAmkilMBXCEk/Ha8VA6QL2CiRL7h/FXMakw+948pq5urvQjgn8xSi+vgp
WX+jFy8AwNZcDiQyGHYhMSNNwyao75/CW/uOwb5b3pBhY4nicEXOO+CDKxdv37ea
v9Xkq6VSx4Gbil2oj8EcO5+KBpi0SqVufgKk2WF7aFOq249rIYVK7PKjXWNcfcxY
KQPMgOkBcf2qKWBYD4OxSCzDCI+wBI0Pw/dbD8nhsVik0iNzWodOGJP0B+Azn6c5
6IZkNm3SH4fMUhluwgMylgRzugFYUpyxntdYe4anVesEO9tZllzILBW/7wvJLa50
/ad3yNmMO+k6ox+uNUS6PaYEYExT+q01drjy4q/i8u3zvM1VtqhrhU5sJrjFmQka
RSZtxQOhcIZeXOYXo/+am6WCnIqVpkUzWT+szSyR9DOIEninFi6w8K6qKAuc7C8P
V/ZPjTGb0bQehuidF4PbGoUBESgI+c4oS3fhK+xqx76tK7hkAZZlvk6j8t+PonKX
Bp4J/VIhK9iZq9yaNZaPMlAYD+1dH5gfqRXswGNhq72ssaLFanjAHJfZYJpDdRwl
EmrEjQfVp1XIX63f9yzmS+Nz2ix/sMu1b++alCqaHcngcqliVZjPOBAR0qQ49rFc
zbMQ1JujaHUEewofwiTC35dz3vaGBXFxqSJfZONL7O/GWsjnki7RYv1bxKxiIiZT
paS3gDHPVzFBaxDUa6dstavm81zX0EzI1n8JN6cE91KmGXLGin0ESDQvgnv4CNtT
h95sU1t6PM7lZgPtTPCx17f0yrmTvF6sP8xbjVh2GafBcdj+S2y9zQButErf3UFr
9NP1Ajrq2EJG//+pSB78lKc5hIQhcTj6K9Adx4oa/8J4GYHFE5fDbDEXoG1JVxXz
J2r5BiOEFDadxH3n750E8qkzEcuR8/2SWiUX2jMg0Fp3/JUbAjT4Gt22uTITf/QH
QnyZbuuIp4aufaFs5GqfdJHnG2XOc4XP9AqdSSa6o8ZAVmuWPopsk1WL3J0NQTYF
Bst/Pq37XRHGmhh9wrpEUqMY2wPp2WxoYnxpT+QyeLoa4Q+iuSdF4Q1AUI0pQnHw
7hMqbU+xgqJTMKiGqWLtQDmrvqVqtzLrP2OicJTQdRCRLRGfGl1YkXkPMyN0HU/7
+2Qcz42r2JjcpwgNDmGOHWOANO28YZgPulYNBTCCO7qwwvQqb2FXEHegRgrTrEbF
sYKyOB1S/YJHa1vwzWi+5VTcn+wXhz/CAlDg7Z60/CG3nUeLG+W2SOq/VciT+pof
Ox+yXaeTBsj1OE/MBPxqpncZ/5QB/ACrRNpPSmYLDYuUlK8JR2rTUcotBxc0USwq
+GiU6VQotznHiqGSRacMKMBQOMmsPD28Xnd/8d6fDpz+dZVIEsvzCDdwtSIEnwNl
V4EDVJW4grUjSWqbZWxG9YlBhUZ80ymj41Py1Ywzbdlsx8QyVSV4iMIxAgMMeTvM
hdeGkAqhlpFtipz0qQNycI+QaT+tgrQUxDHXwRFNCsZ+txGdvqTl8rZSzeO0MDbC
LhYIj/dR74uPbSi4LeAlzRwjxsuwyYfnIfhmlfItX3mHgYilzuxYZL4ZujF1POeH
cuUQ4HHhqHmkgIRpJ36870rBHO/25mQdi/Oe19ik+1J+bX1lmP01zfjJg0LTedQM
HnsOzZTz5xH0RAcmciI7Y/OF+y3pne0PtV5osrYam+mBQFdGhjZwFwjeT3wGioUK
i9vCMFgeaccxhfR3mdA2ic7834hD3R+MBHTgzmDFSOSr+K4hAyliBWR6AS1eqmtj
I8d4l6ZM/VTrYKxSqF7q/PBJO8UNbFcu7I8wOtca39lwnnPlzvzcw9phPuXfyE9b
59DDsOk5YjtNSalo9w4BRlgzBHrQehMjnBrvZhkh+o9Znj1iqpoIUzcFRdFf6yWW
mkDBvH323y6/OFSNujnPx47Yowful9kQdyYLqXOTHLBezOKO59Z3mzLXst0ZEhcv
UDRmmQQ+r6yzoGoqy9v9pBFuSLA4JkGxb3l5FznBqN4ieF5VSzKx6JV5zQxpXtkp
oAOlyHyH6xtkNxAtx3r3YtDqBNfAbLz8j6WkUod9D65gPZERqKjdbldM3OMBACUa
7KRBikoq3CnpM36R2wjVdn6TmwTpcwBgHUwIrshl8shTTxTYJ1+2yGydfSx9GDeO
7LKfZ5irsqAGs6HNmGLdxbuDWm0cDVXWup38iGpQzkqZ6JPJ0X8IaR/19dMlB4Ke
P31DgBiietCdv7ygx6nQ3rfT4kA4Kc6+UfgEWFa73M+PGOjwuBXj2vOBEC7B6+b9
a3VmEiOF2eED9Sgmw2gkGP/h2Mium9Svo8rg8jXytF1zeRxOnczPPeo+lpyxvnu8
EQa1JwZLBoghwm/XS/pueVN9MOwUO51p+9fLziYur+8IqoNvmwB3/+VepNyOrXio
b1C8p3n4tpbo/TwRePcFPxjkdwLHVkV6af9oLe8zkrXgX3+3FMe2ap70DAjcMOv9
ejoEn15+hhb82bDDhAou0bD2BrkGUUU0K8SzqVA/4/t0v0UQNEoHwsmS3JrBUUdo
oWg2qes7h2bPWnNilJA5cVD08K5e4erP1tyEKmOUGYnAfMtzryU436guxLcxqu1j
dZzEfidQ32Nnzig+XnP9p6uCbLUVBdEEYccWeEg21Lm/qSrttkb1IvP702mW2wTo
oOCaiXOuEfLLuLq65+QD47yCABITCxbefr+TTsmcqodVGzxnyJpz02m7vUpDLDby
IBWsQ14ME8+ve+95tYiy/l/RA/em4q3Y9ImY+gDs4DvzSdkdTEP0imFdgRypQTT7
Fa3AkalQpCzSZNDfJZfHW6wdYB0qOYcJs0h6cWdR43DWN2clE9AbQzrM75svMKh/
Y/1NjqkLCERjanSKYEBYi0GLpIgZhX2KF8RakTZws27NLpoqiwIg9DaSOXZnvbWg
20+pg2dteogJKABGRlugq9vuxdziYfAYKIiZS7FYRky2CN4WUknjeSzmMYj2vtxk
vsPnPFE5pc8+fykC4pxD9P23mhMpZeYkw4huKw2zbIYEWPTbwjkqTM3iI8+yxhbR
xnAWaaZewkosQ0kTaoJRE9t598qP8eFUC71SW6gXA7kWpTiE0p08bhX+ryeWG1CB
MwvkSn+KM/vd8qTsJKKC9Yj+6UJQC8wjTev+kQ+qXfLg04fecaNzpvF2/dX3BBxJ
yKozBbekVMEkTwGGAhVrvFCY4C+5PCpcy9gEZKO7fD8Bh2dAYfDBhW+L5vtbkCMk
BPDEVrMif0XnaDmZo8V752JQY7+Riai/Z5Rj+YuHuTd4KRetgtGyGUTw0U6Uz9dc
8SMSlGHS78BZHbTOP7zwVzaKjK8By+uyLjwLEux5/BrtX/0IeA4f2fbUEuTTctvY
7w5RviOsauzcE4bJH3I8+hrRwSP24VkRtEay1iBqlowxQmRSWTw42bcAD9p1YQoF
tn9nEbUtnmKz6Rh53wZP6B6hQGxQW+fVo7RR0vpSI14JuSkVDppevJKsZWkoeJbZ
ORgbuLRZkrLf6jEA3qVxRPwGWMe5i0xtWy9X/65MsM8KFVoTl4JPBrg2LdfGjFFr
xhljC5qAZ3ANh8FcNUARtSib+wpojfOKnbDmP8dX1vhD/ytiudY/b7dG4CcNxeBR
1mSBfT6e0KJUDRJYVWSXto5bxjGIayBmxv7z+tRJOR3xEdSvx8kESXJC9D4O7TW+
8n6l8kBKpm0dP1fC2cmwWTzkaVa2mzOBS6NCGsy96SL7Cj1ons5DodR7DOmz3XhC
LzqJZ53IGOfchOCqoZgCUv2wzd7Fvv47xFq6MDMKX4WZC2dc9DY3pcWB2GqGfrjN
PWAW1HZzRzdrBVbF+Jk1wpAwmEH5wJF6e2bGj/w43F8f0L/HZwlIZdbW3QKVyTVC
T/5DiTHqSO1aetmdUBAdND88c+F/J5GbFKhVp1Rc7oQfIYwWhOo/cexIJydhyoVG
1NE+NF7cFExdB7vVRjrp4phkUHyxxACgD78pXYiWtLDonGiVYFry1s71TlId8lF0
DLHlJb2ZZ+QHl6m0hcrCWFLGxtAS2fQkaaLFPeLcs8cI5Qh63Cz1UzyZJ/xG/cDF
F6vPwwjTbDWHrpArjdqrNQj0ziq0dMjT/kFtT9mPevGmN7kaxRhs6sT1M9o+XNeL
cnH9woVBBc5euky2WlqRPS7vTHWgEh/ClryUIr0PMHCvq8NyAJUqlMEoozbZbxWA
hZg9uxJ6gX+1ZHjEbVUyBZ6Y+1ShL+T94jfagMTVEEJ1A+3u9Q1bdcX/vRiU/wy7
tww3jEu/wADENtYOQ70fDfjpLM5Bp9doptaITdponJ/8gqwKB2nMCyVCOf79oz2P
mPSQWvljFvaszYkwWSBQ8AR9zr8FhiTKuSrK5zig7Bah3ycx+5cptXSmUnS6gdie
afjyp0TZYsD+RR9nDNbNWu92x8LB4HyCMNthOsHTrE+v7nfWHZoGGblsRxy64iBa
RftFfQHs7jH+K4qH0k7/sdEixWPvWoeGDVa5+WJuLrdhu9VwKEfTfhPxhU+Mjl1j
y+lqQMESFsi3WglCNAcs39SXXFnrrZ2AL2Fn8jLFIm5MTKtIAw6PLZWT3nm/U3G3
pN4/y3SXWMA+u2R1hCakvMxc3Rv7tbNIg9jYtd8gBU32kLWAHdocPdw9KCpYtcHK
PynAuP6bVf6S7aE8Ao4ZUY4WIi9rfGTsjYdyTJI6Id20yQDElGIyFvNAjYXEIukr
/wEtIjhBSFbdzYBtxMKdtDRT+fwpB9sKyBA+RLzpxyFkOskfzYPeIyrpwq/mnevp
zKTt12df/LkKLpSsMyR4asSJxSzXWkm6kg+96dEOJ31+QpKigP4pkBxjgtxfVwf0
DAJcpMYVuvQkAs1QQjPeSOLu+SF7FTJjdIzcd9/HLlrAmZezUwugaYY9mTw41ngP
aQ2pajz2BMjGAqXKC3w4MUQnawBVF2Zqo6SGRKS6Q3KftsZMcGbD1zokqIvGWoE1
GgyqrmBJTLPgm1V1kwjLYRLKbu6OKLz66E3G/y8lp5MqR1ccvDjt4dZ9FR2h9axR
TUMrLzL4ozGvLak/Fk1fxzB1I2gK6HU5fUMxj/ZvjutHBiWkoTjF7kgVy22VyoBK
kx1USnjxconYYbzkfy4wHQ/brZHQiLOvbVwp4PkO7hjY4ZRIFiwfGw2BckUFUwiY
Mb/Mtyx9pekrvJX+S7KZXLQjA5pB/jrKFCtyvwzy9Tif2EkAOTJYNySGOILukc6w
QZMqS2E0StqdH88EsQ2CYBVy3tvUvvHyOoe3vKSL2VtU0dhB7sTY5VokZ2uoFZvi
VFkDdfXZZnClmdS36tEE8FzJvCkTkFlCLvGQwpPyTP5SmnNLm+yQ4KpLEKSeAaL4
H9Emeq2zCPL561u3xwL8L9H9ChtGagxZxrJEC6zeZuI4VqsgdJc06E6vKyxj8tl8
vkSCztHht7JWp8vkgJdQTvuy/1/uuv2GL2athVaxqitRa3DJpTtjs5LpQ7jGS2rj
RhQcjKO1s4pE/8q6y2zTNsMQ4Ce7NVUdA3TQ8zIm+W/QpQb6/jQNXjU2tcO42ux0
kkHBoFaX/sdYXojCM1tWAB9KcPerFa6vNcvJFDorLTb/Qlzx5FkBvUz+rWxVaYzc
rIKoHyQGX/tO4Tuyp+jLcm/QKobFnvereIoWnJWG5rxHTQYnWAVdZfMXFamHx2Mk
ImErgcJWNyQgNcRJmRSK+aUeHP8ZUDwMKNPHjFiQ14nN2ZnbU9iz+8K/VOFYY08M
jrG6pXjpmptPdAKp+QT6UFJrR1IK+We6Dyr92TCTOOYm1UEb2tHayE9Ayz5rLruW
qwKs2b6n2zhNAPJ/5uvosinnabPPy83qKh6mCA88ZTPdG3yV6H9HOGSZxjBj2T+M
rpuxJGdAyntPM6FdmzmGTblEr/bhyFijdgakdUtNiGCJlUacr+yIDLmspaFMHhZf
kyH3Q0OzQukaGFETgT9Kk8VClnNZe04EPoLWKlEG1RAUd+Vv2zK9V4OzskWuPuAC
SLM7JNFqEMKDyY0P0VyADe3ISOaTlivJ69MKP8US1vRMViUXWUjobrxetOKQiMqo
xP/l8N3Q8LNJ8ruv8jaFZCaxl+UL8XgH8sTeFgZvBGXliZVD90Dhu81lPBTO1jRC
siHS3nKFIGyX7Ff++MpzXxx1RPrq0kPk2YLBr+gyoCm1Iu9bibk+uMHkTKDHCUfZ
QtTNizMYX21t5kEQKO8ni0GWvpQf53PPkB7CEv0Au1hd5FigszWbBpNTpGzVNfRH
5wbUvoCa0bF/dNILMJPlq2q+CK4Pywcsdz22mLnB9SURuz5CiyCIapHZBB/XOR8M
MioYbACQ1TkwlZOEg/ECdGHbHPS4Lz6LvMYYVrPW6fyuIxkRwzkZOPkgCbi+D+rx
Qzx8UFSIn3Mrhnf58hja5Pb13BkgyAV0xaPknHV6ArhvvMrFZFpSwMNJk/AZfqvg
5ucN/tQ037OPiUOtI2rPuDo+w/6EDFiCpuBjrt+qF2pOrS62Jl2H+sTYgru02NhA
vg5hYGEqOiSxZHaGRFKGVcGBxi3ok1jgmF6bJlcXxf2KtBfCvQrjl2t0NH16ECAO
gDps6GAzVFiGzgSTl25VgZN8gKGOyg3FW9h20Edwm2P/0zTmD+zLCzXZ415DLJ2j
lUw3+7uADA4yXaUF1YrR5SSjpRyv9s9kFm6bwA+FXR2bI/4eA8Bu1ksAB0d3qD25
MLfREBCu3fZU5OEDnuMWKAQ5y8mbS2IQkR641zLCxeMgKxNxvbBeTbXzNpwposCM
ai417cl2rSn05CqJ9ebezUYzOve0EMd6oMjeYFwpHLFTZnUtJLpkMf0hxC1S2uDk
M8WhM5h4xNyH7PK8iNhkLrYbnkQHTMm4yj348GXpmIsKuFLi7ejbPu15xTjIhNkv
slrNg7fcyTTxsaQUaQIEkwM9vkmudXErXc7DXeL5stmrTTeqApqfupfpGf3AVUci
Hp59ohQHC8/mUdxJxEG2kGxhtldGT4ZrD71A7I6O+5CYP3vhSlkpOwa9IVPcxyDI
nCK20xWXbCzrwKlqPekHxLFzbGecc2kJpJuVzZ3lnqQShV1lR/AbAQRL6OdflvgB
PVgp/kns7OEEco7ICZTS3r7crmPsJt+p/BmQm9WE5/+85v7hd4WiTWlo3xorb7kR
F1Yt9jClM2oTnHTxnlV0KQgJa1hzVk/tI9driLR1fh3VQJM+n4GKAxZ17tsBtGcj
/yPYkxsjn4dzXwpn/W59GqBPBziDWAZMa19Dbp/WgoPdfM1KlYf5J4IWMm1+T6fk
1M6WrXueIMz3A7s8IZod5BD+fvcmZQ/SfZegbma0xFyCjkAskDDF6pfSrt7l8vIN
XUi89NXAq+nKXi+zrIpWc5ypc6ACKXy+Q50TvudlSLjl413HHqvj2lxDdMk6dX5X
b9FJkTdm0CM702k4f8/sr5DEDPWhliarSu/FGVk5S971OdF+zLJZgMqP1mp8vSjZ
WqhFjvtfV+KprLa0VVNEYQ/gEJBvaSHXxVOosjR9Kyu6RYAdStKPXWXTH7WWSe9k
QvGbzTswTBDQkISrqSeWt9fbycYW3pia5r70BxF9JEv2UpCVYMzHpaYQ3spSEFwV
We571afAwiZtlPBK2Z0PJD91mTAluUEvLQ11YSXKX5a2sJtaFN7gpnB9Uogva17E
PUWxUtnBgoBdXCtLvhROLx8RjfLMo0GwKLygvMDCzZGLDmnd0zr98b+FDaPTlnHw
YZ47q125NqFj2LAb3NJKaSA4sXPgaU2y6FPdlLYZ0PfZhG+g8oJyA2tMPW1gTiqA
0wE9DbvTSaYQ3SS+LaWUJneEVSNRE+Bjjtp+HIkcCmfbTGVaKO/ongWy9bHtRLqY
90YM4fNKpOCUUlRPm+VgpXFeJw1eTjCYCyUFeG3387envqSYQ7ZNwZMRgg2rh10M
EY+ZRsxS4hCEpe9pdEDJZGF5s9EYP3IgI36/hpeEO6sZcbQxjW6vimuKb5lirMv+
vFMF9QTjbYf7MwL91t8MRc1ytJ9BnXi3WcSopWOI+xmwBgInlXtEq+DNCMK2SZNi
83LX/+WM25m1co49Qdc+uY8bn3Xpe/lWDxS+wLuRGO3xlI11gP6NyPDlaAsoMk2j
Co4FwbiZrAdXCJZ2zos2GjjtbF23UFRFS7dBue9PMeqpCwnJKklSSgUxJqTaK7rk
7Vkf0G9ZkWxy3Z+iI9amQYNZeLUin+sd+f8YyGJYqe2D+uqjsY/TdR7bSsf1dc4x
GyGZ6T2UI/tAwX5GGZwhRc6eMuLvviJHhcgilGdfj5uFxUxo02fHxEowm+2cWQY2
ykhNcEXTFGXQsO/P0WfIhmPNfb1nsp9nG3krAugNqakxLprSM2MvAkvMKJWfy6hq
CR61iyKzfxiG2GqNy2cl8rzv9qECMDrrLrGeQ6vlMvLSaUN64EHTx7JSOnsvLUPp
ZEytU9Hw/l8PadVVFO5ZQ6vTckZ+JLsPA4iR/3aNTEjuKg55RKVQCBevon3N2Z8a
JVp//Ki0gFIYeY5kioq93mO6/6Xo33fuOugsH5sGi3sT7n31s1/SHOxI3seyxq40
SHOUUysNiZTe4tboNqLxqpK1HY1wmubr3YIGjAQHH9t/TCSQeKYJw+t3rJcO1fSz
CTIFhdUB1DYn/DOJ81NaZ6wptl1goZfnwJNqlkYS3j1/ztFgP12Ko55k8P3x+5j7
ZlydU1tpAyyTA11vT9KKbySMhp2SiwXEELISraI6Y4S6/kPurjpdswRChwIkN2dO
nDtmRHDqkVv5m6kDhX4kBh1I/P6yRL0QmXXzfu7eKcdO3oH0XquydqqdjSlt6WZH
4JRis2HpWFHTdmx6eIZVW9b+1HklTc/9ETYjsajk+IDy5CyJTCegSbN6qU0sWRsc
5eZ7yjnZUeG9ZykXLrlp2NOtQ4u6OopUZtKjCqmt4CX/nngm2KAbEmk4VUjIEbxy
8HqKg4r/P9RSmAkcAVsrdCtRbbKt10/AC7wMztdSnNwPCe+EygzCXweoQ9+6dmZn
Kzc4mHNl9bOax+0a/PIqZ/vEOqDV55Rxq50hfxI3vphYBRdRlFI4ogpv9iXs28Rv
LtCLPCgIa2Q4X5ZvG35rRkwDTb4OJN0k48NH3U0U8OD8rh3ArAPat5pgZLReAxRx
q8zqJOwm9gJ9SHK2m4bY3PHWZJgBfBNX1E3/ZtT6Ljjbov3zZH7102PsI83DkLju
d/3qRTWzutiVaVP995et0bRSqG7Zca/9qkZEC9NlnlYFgJVutdvs46yFPy9hA/uw
ReHHWGoe5gaiXMst5/TshKCEduE2gbBVJF2Rsw8ten+VWLkaZadpqKpf3eXSQHYn
VJ9ukvGPrMoq5ncRaEkhlHJwlTW4VWYesDvz5w8b0z9nnS1ZGH47vdPhoeb3+m/v
4oTa6fok43qVhENm02PSb9Bp9ZhsJ8agIl2HceqMf7ij2stD7Xrhg74nVIsfzXBx
GxLxI/7p1I/KhlCX8d4u3I6kCHFyuUwbt30G80QwgpQwoTpM8Edm992ww7agB8S4
2NkNhSwiuIGPjj1MNwTJOFOzyNe9/J+3mJmx/TFSnXdcTBrcJmiJ3M5rp2xqC1Nu
8C+NL19/5tuL/GcU3UAYD/mhe3mvSkj+r4WpFAA+ClquiLYfwE/KFS7YMA7x10xJ
4AGHyQCuzl8efvlQIsU6wS71NFKPng/l663k0potE++yKzk8HhStkp8e8JfzEnu5
uhZ+lAJaaNTpTnuJxupAQ6XIj/DHGEL9dPJn03mSOTNsw2I0u9bZBERnUR39FzJM
uFgCfLUsZBzkfdToKmWPakscpyb3Ybr9D/8DLTdhdXmhZsyzkrmDDhdmGE8lYJ5t
XRzmkQbMHOCaOaaM/QvwOI+Wpvy4Bshm5LbxweSejS7patdxWGEI75holClY9UWq
3/B3mYkQpPA7PrpJNJxsKEVPfQOavc49Un1d0jaiqKFVNq9ATiE/HB3cweTZOkDq
vPIp7GFLtl9t9hPiYx8c3GolByoD+P6QtyXUqTAVZOODqZygFx/wNYxW1yG6RNkm
aFXtC4nLvaBnpzsymlCQTrwa1PbQOrssP/bxaXy/0zwRLZN8CjVx+K0nolSnfkJU
utLEPFx7LoMQhEUjezk+NmrouMSW3CBMteoFk8CCycXLiezyiRzPcU1B4HFJ2tSS
h2GAZQp6r3Ara+I8nO1Y21D9dR9DP7rhK3jcwB6AafGtsEAQpNg3NUtKj7Tvo6rB
ElEJ6Pl7DZKvef4fmCvL6WiL4bmBbimUVvRESpJfaPfPAWK/nASU8C+npuQAQvcC
tyDp/Zr1KWf9g9VWb+I92s74dB4Q9Fo97siQYF8frc1ppjPxSsVxhpSDnbRN1UoD
S+wZW7gBwKgBBjc3oXeg7N3mOxG41+c1Jh8zgzsnvgd6v9TP9WGQNq3lqpO5Rgt/
FNKCvIoQJ/cT2MOogZjhRGnAFMwmW1UnCsRFZ9gsVWZjSW1Tpf35mCKo6m6ckW6c
WIGKGXBg8glRI/0wjh8UQawwjXdV0WsmabIgYkFul3yaOWUG8I29fFxnDrBZ9TK9
hh8xtS7sBYQhGlEPonf/LiWz6yHIGDN8QQY+JRHJInFXpSaQh9cQvtpRAoe3h5bp
wjbW4jxXypRTEP30CLKyoagKWlB54ZLOAJZasa8/C/fPj5OPx3lTsoIOo5BS2mQm
8JlSMQnR4hV6wheaxaKVxnh99kZa5Ze3KZxtwl9jmTv6DkFeeAw9TBnpt6VRS0+U
OykAJ7sC6KWlEB3/FPGFr3xUV7goCppVWTNSe2kNI1INcUIp2NuZtvq0sxpbf897
PTUIM8+2rFsuZnbK0ZyUmU+fbBs1QYh5hVlzAShV/1TVj2vRjCbq7vBK1FQuZI3m
kqj5xD2jHXkd8gRacmFFrdKQImfBcgeYC2Z2kc+EaDpPw7epSFpKH+Gg5dIJ1Hid
MqHKvqx4aEW9lxBXY7XAda258xJ+OXAYI6r7mMzeCqzkpQkQFEpZ1rJTneP5U6+Q
Bg+4cqLD0LqLy7sLRzwhgFvg1y0a15FoD3gY+Wp822DhevV9GQWuBYasHbU4MVNA
cjPCKoCUSd2l/m2NYJct+lvv+C0cWci2vGsl1pkzUZ77i4zQbEv0uMHyTzhvN0bA
TJS9F1vyuQhaMDSw6RhRFUTQ3KdmsjWFBuReoUxourNlEV7CVyK50aVFU4vMsQpx
hGWNtkTJIVj+vT19sTEbtzOfLLp43SOjk4RVbSH6Yg3HO6habFcKeBIQIhBTo/ZY
2bph1RdTHS+puFHE+2Jx6CS1LUVPIxNIEGQb9VNkxOflawyj7hGTNsJK6MTO5gl3
5yF72lpOzueW7CS643u5mOEe8cLCgiLXrR6NCQbAijj3FaTu5a1EnS3E0xL6F6/W
S85Z1ORG29UnV1O2oHECO/VnTyH7T8cBLEtP3BSspe4t5XSKZsTL/AB+GJkR9Z6O
DQphKlMibUEEcPAGfrciVGlZ8oyYepar9cRNRvDhEDJEbN6Q5n4kQAJvKXjhesWr
T6y7deGof9A8VLgL3h9o0zhbOziLsU07wZ9Y6E9tcR2dMwGTCEdnAqUdRwnDB7tm
31wL2DGNO9DgpQdjqY3WkS35LTtyUO/WKsk86kGrqZ5+yl6OiPZEZhE6cHDTV+ox
ketoHOyymHFujhXTWRijGX+YIzkqtNmw9ZhfP3Lv9Bsb2/7RTYME/8XThiIPbUUt
Xobu1g5Ibc8tyoIYDzWZgiGLS/0XG2DZoya4kAJlx8iXt/lTFer1+juoYgAZY4Zd
H2WMja6UEgFd3Kh6tGijipUIDs50QM+MMkGU+SJDAXnXVfILbBx+u78z/DpHU/W8
yL7V1O+9qbCsTH0aF7Uz3whIfL26TRpTFgncvodbA/WS7RTO+SOX9vTiOGxsZO2Z
Sk0iEk40K1piCM2F1QFvz5ArydUqh+bRaPxiVh9KAy8r3R++NTmh3YOdgTH1S50R
9+l7Lf68E1QshNr9g3si49lhlk5/n+mUVHy+PYWpaVuNy7gYdGIQ5Jcb3l4A0bAQ
PRlfpPMbN4O6mWjDsRIxQAjhYyyX3GGZBa9lzWPcip19xiQ/KoAcYX8Z7BG75V6z
HlIKBm80ZcrZS9PCULtc8cRx9A34LYQ5mbl/DA98haOQkuByFOU2EYYfEs5PTz9X
w/4ZNYEGgu4CphbQYIidsEbJ96gSk+ToiePbq9T2yTtq63yeRkKT8Uj5Tc5fxZwH
Y8f6HpVaocImXawF9CKAoyo49LSOJLUZY/mDle0kURL9k576eLEqpD2lF6YSYl+F
4IirgRIedG1Srq54lFSSotJbPpQOWUKXiv4NoJf7Spqzpe/jQAepFxQ/nsez8Omr
P3IZ9AwByP4EJSBj2lHXKWL9xT4Sc1cJT4e3Bt5J32YVUWkZaOFp/lA++wopl7XT
csjetjMRdkgOwrQ4cJ0fmvM65gvCJIev6LM65lOBPFpOIn6SJgMpzb3zPodbwx6w
FTmyPslJFMi8ZzpnfSrkz5PFfu4L5JQWfSJ4j3f0DN6S+u2YkxkfztKbKFg2kotn
ftotlFHo4TsyQ9XUmtvThia3S4kmD89y/OEcQzagOtvX3xbreX0Jgyuqevtebzv+
oWxkDHlHTqCuhpaK+paeibsfl6GdUsWGtbg9QOU9/A2bJUOeWTFdcsGnvA57S7I7
jNuIHdT+Xow6goV0moVOB8YU/CPGaD0YCILHBrEhSLfJIahj6jvZqFzXo398jmlt
fDk6WuurSkrvm6jk0tPcK5E8cWVkYKknRuCratrSZVdxGYIjUd+d8VFUk6pkh280
vfUmndJbiyhZa9MM+97H4iwlbkeCTfX0kpd2ZnXE4VCGAd9Op75ilMxm9ldWmFhI
fsFYuhjtvWvX0F7Ze2X29vfCSlZWoMyIH72uieuA3RxSjEdbmSuJ1+qUqUwvv/Mo
oTVUiBZQDHwNHjZOOM2m9y1dfGKBQEparWJGeNXe8iRBjEreSZI3a5gVXlHIF4u0
co6NtQ/WuC7rXP2/67n3GguQHUGO4sknu5WGuLEN999kRz1x7JATjUesJfBWr20L
1vvfp+1Vk/kdbV60idUZfKtmmUDg0haJ29MLmNYR2VJGq0p6QxnferV0eX1S1W+r
wK8adPH9cRCWYgnluZrJvv45ulv5j1x5IhoDLVcNexyQ0Hr6fz4l6mf7gV4Wfp51
/kF38q+OaPMbkLdvjw/dNGa3ps09Zcu5DPUSnRHknYRySBbnwbzGsM9Q6Xjg1eOn
CgB5zEcobuoyImM0NWS+ALbLgfBjQs53/+V4t5+MbNA5+mx95Tv4MPLmfl52oSz5
KY9CwF+IPoj3S8FOn3vIVYExkomqPC3PstkRZivZ4b2DEMQX8KRVJ3Pc6FgD2G/f
JI0S3VnZYhed0kUfkVhEMjiabU2OGEcZMB1GhDtgiK0XlOAYnjzvXpIMSOhy0ihs
kZ/K3XzqWTt9El0Bdy2njXtb9Howb21s8JNgb5w1jFkbTfmbOfGNerOjNVa2r9aD
2yqnGHG2CRj/YarxQ0R4sAfM4sep9YEvmW5oKYQC/mm87vuBGi+vrZXbx5WrrH1x
l5EYcw79xcXPgI38CumKpA3TzcqnpaXQAtt/XlhGla6fn/oASCOUOthUJp0M3QMt
/5SiQSZaLIm2Y8uRz5cWsl5MHOISFmrZ91PkOdrWxHnYHIFpUjOCj+hMrUQ9Ye7I
9ONVEVP87g2qtS7y6nLS5ujrisIdTp2kSUJFjjocfdW7krsPUYr0FV08pajHMWzO
i8eIUTlhrEdM4TiWj3BvaRLJE0ZF7mWMiqNyzmr+2uaUdml+mRE5fGRtECtIfzy2
BXzNrCxw10ceDEZRSEjuVkk1RwoY8CzGiHL4mqo5BTtRFpL8WBJgIqQdp8DAHWK+
1jnv1hX9L//qK240cOuVGzW8HUg62ha9zADAelI9EDcj/YpyhfZZXs9NtSpeNF/Z
mxBMOg2Usvc+wHG0+D3cSC6URoyPymaM5hPO262RBdcdeSQadQF02+Ega6J/hx8P
t/s1HxjyxalcRs6QpkWelljDtIzlmQ6j5koA8xc6Dz16OCB2UG52GaZXN3wwaxqN
5x8jd2HfCJO1pJ0ROf5p7xr/LN318MfoQg1PjbBnMy+gdt2lshnx1L2JMw44dLLt
rLD4KOc003hd+TaqwbzVu31oiUuVXDqMIlLAGG/jYVXoCHn40FWlJ7w/vVs/KoeP
cuAMXEd33bLsxKVP90WYvlNJ7Z+P+sQoCGDyxWYPpI8wV/9/sDDiaFDv4rYNVkGY
FO0uIuQeWEhjt8a7G4hpAWzeYjbvYsFo/zGV4Ex7+sN+7Wuk3ZBdSwWpu1Bld+cN
lmHa/vaO7H9aiUUEqVPzevO6DVYzRREkcAeR+6OhUTy9DDqOiOPx8nJzaYQloTAj
NGxbNr8uPNM2l2jkrleQvu3iqj19wJsx/EtL3TWCwfLnXQ7Mfch4GdW14ictNjen
5MotgmNhgjgEjIRgUkbBKHLwnXER3EbK5tcNHnKopnfideTLIm9QrjaKMof4x6Gu
0MQ+wBcfmndH4AG8TvUNdBOrebbCppVRE/djVY4k/HwpQD7SUmkFIhU0hixD9ZjK
vmySxK41PMLLlMRh90C6ClqauV3fphCf4bDAsxPYN7L3X4camhsP8I+6L24gQcPI
/KKz3EYPRtdYSEzdhX2jBvaafeD4cosB6mr3Qi+MLon10vV5LrB8T0bRe6Z2JpAV
4SEd6JPy3Wu62jAvtjNiy+do1ZNX7Qwh/l2ZP7NEOePBUQELJ1VifdmQl2Uztq64
hs5ZTlo+qHEzwCOVsuU8gLnGb0ti9PhAdKE65/ZNj9DFaScfU38larVOmEi6S/PZ
2V9DOaDXcrlaeyyZGqJsXwmR1kYqzrqkMspjK1qnSBV807i7OwEE6UhN2WoVgO6B
d7gy6Z6SjUe4eCCbQfhqkFNJ13FMPt85bBKJbIsjeTgDjkeimBotHr6uZ0Yyb7OJ
QR3AvDwuQg8yz+zESovhTNARXYZtOjCYk5tAq23BLKKV+qizs9CfYUxL5hNeZiXs
yRsNTgOLBiPM0Ji9Jqpbo0cfsfWbXqtHHgEecyxmVD0SAmSNNobeWqd6uKFFsN48
ZhpqCXFuLtosoVh8cSfPLgR8gdHAsKgmNMUnSDz61qweKGCyzpQfdM8VgimzIQ+Q
6ICxgd8d+t3EmwX65VTWM3YK4knctMa/292tEM8MJZfKwv8pXNmmKzG3+P+liybm
DWDpMKF8rzhIfMoF8+n8305fGmZJacRLfBGaNApA2MB0iR0u9sFDjUC8i9ScTmqR
r8VFch3K3V+K5hV4uTpdpVLVoY53C6ewzjE3D/G/fEUCzD2zOPqfyGriYjxqiZSi
C/sN9dO+BqnUiu2pNotRdO7StTiQfi5YQY802DLZysAShC1WBZviVqMDAj5l4onc
QECa7UG4OuGkx3NuVx9gDxQmRf0g0WgtDgwLDsFq3ZKtmOw/51cHMImhDBz9gmtL
i0pDaG9n0rn1c/ZJgscj+zVkABiN/bjIb6db4IDnUgxWGj3CL1bnYwUiCnPhbzsi
qKP0bETgsLUHRWf3OVQCbR9zk+cUfY2RDUyNjJY3cuhDdL5KuMYBD+gklvg+iBCc
6+IU2sP2O1W3EhgEQCD0WARpu2JVAylrVqMCqqfj5/xtfXMaLWwEVTBAHIV3Ecjk
YZhgXIJtvML2oFkrI3saw7QPvEA8EPu+L4CTGrAQc7cibNHO6PcLvDbF4bEnIShy
7OUbS/ScZ9r44OgVmhvvhHLcydNGByi/nbAAv/fb0YU4B5lTVYFGx+iHumO8rWUH
LE50wB4AI4RkLHYU3874Syzk5CwBoYYnT7H0PL/GEawWt4dwRITBKeA4oAWtPXOO
gDYm5M9iyzVtDKnc8jACIV5sOYdysf9LltQv/Z//R6P3YnTskQWtTe8QNey+cO0V
Q0kpTtN/ZIjJTwidA3lERD9FqvKGhXjDp2bXlgzwp+0Zw4JekTMyQw1plfifcwnp
8nz8iScQtngKnhLisE8rhpFMicOm6sGYLA2uwzT1lrcaLpG57RhhyoGiTk5Upley
0Nlyq1dZn9oXXEZaXr7uecy1RaFqMnUlFF7sF0UCCOHEspHSsKhmgjes48eedVu7
TpD9W1qWPDLlnwMoxXqS31jCIyuAyo7F6nCXW2ES8BdaJ8AFWzfcbNFHxWrSNqL/
+2gjv2Sghx9O8Tcb1Uk9we7J4IjjqkD1toFBZ+4d6koiwpKC/Q0+Scsz/zRDCV2E
EwyoW4jvYJIh6hl0hU0lpYh9pcmwkyD0nHNcpNtFaFI5m6R56WbR1RvKDfJb8BuV
8FDoU40SU9GMK7XGHe9uH1hynRuMCLZT5Q4YslcCDl+3XEy7lr2HfbPHK27NyUxe
7xWOikq74FRs99P8ChxvAPoXD2ahg+fCEdIKRuyPTe1SCqZergUrp30YkhqEIsxv
MZCVXCHXcjoyeD9TtmH8C1w17al6AjSUPOdKl7v4zYFxKLtD+St5vLog+4zZFHe2
Du1yoMxzKkD0FG6DSnijUt9w5g95vbdjFyZIfpG2IMAXS0GbHbuq3Ed6fl5U71ot
T2q3XgWVqMoqBZPVR9tDYYSc4ZtbTM7nvKfqy9m7Hk1TM6MvbGijB0LALF54W9He
d56lxWg4dViWkL11lRENumAtnmYuMDu047bDyP3CM9hbcC3bw9QQSNNdaeUcMASQ
2WJYbGcx2sM8Pvb3+JbhW/Cd9epOYx/oerFOSNf6ZHffiPZKnXrixmq9NuDdGzkq
qdqaCrL+C/1NquQwPX4qj9jCmBzlkuTfqJoXRXIQ3SKEVFrrrmOJA6pJx4NBeZ4a
ySkkXz2Fs/9bUu5MHZWyEbtoLRwRYE1WTYFu2GLWlW7hN6SiigtxtEherk9WVcIZ
Cso8Lf1WtJeh2VSFwvSpJH2ZFbLaYEPByV2xPwltMcmnXbd1uJclrYRLZfHoGoFy
0XqYKLWJOJ7Xj44SUaeNMAjGVWD5mOU3OqAxtFKga5kl0GcF6/Vb9Abm39WH2H02
f8thyk3OIwpzxO3SS4S60PP31sBb2Ykx0uQ35vmW+vWvcJ6X+xfRuzngN0pnidPH
fWsR1JoUk0beXaR/4g0OSzIaqagJzm4zpVhdvcfU7zzsjT/B9SXIzsrSJUWSDH9V
vaJpMPr6wxqQxgy3Kgm5+/c0GIHAUQ7+Trv0Sz5CM1kmcHlDDijWPKbp2wF9HMqF
mDxCdIQAbimObXhDKNEc+Kf8+DQ2Qe45Zhx3svILaby+PDcR0ku9s7poUqIjMQtJ
PHaYjBCOX30mLiH4oAqDPrV2Wlp3zOMgw+0/dIwkMfaLYcj9E1Nyiujo3I7ZekVq
qugPFwjzdSFrE6TPzQkTqzGaVxf7Y54GB3at6O+/uLdYD1XeIqbyCMCi398Q8zmL
KC7xO/uCN6+Y6ZTccea6qFytthKk/71z5OEXDGGu+t5ziXNgRjhEZB1/ribti3L3
KLRtL6wWIzSaCAdtj8cHsLB6PLz3AbJAZasDZMeSLbYHbrqqyCkUitWEMhwITIDG
axJIU7w5elS3PsFbVi5WbIh0w5RlFfvKtHfiR2F28aaDQDNGR0nFomkJZ9wYLygd
JCEDEJwyPHdQygZ/sdVOBMkXhV6R57Zp5xx+kMYZqfNZIX1TYZr35mCn6ocpX55w
t9OX9Njn3g2ZT+GmE0yPMnT4LYaqneR3sWcZk1Di5hO9FNXzFVNAnaRPcodxXEq/
Kks2/cZ3xwJJJG5Ve6rxmnBVGRUak5hQZNKxJyY8fbSOCiD1XKrq2G/C0MTTn4u0
m5c7EvPwXmsaudoclv/QYapDaZ0zvXdoHUOadIv3t+ZcoJ4oU4D2fzmGT8OjHgjI
iOtR18EKMmhXWzCuf4emBTP4FDqxqlGLzPIgw4llYnw03lxvVGZubIVUMEfP0VIm
mJ1Cmh0jWiDNqEhpaNMkywD6pO9VyysfwgoPPRsBVmdq5cTLmNCagwvo1OAD8moC
hxwEIbsUXUkUKiKQAqNq7Z4sL0d/eW13t77eGIxvbe48QPvTJHvM/2HUrKh7+qbo
/Q91LeL9m/V5huC1bCJjJfwHI3lpgCNfdip1wkYRkJBJJNwmU79KGKwTeOezrQUW
QHUGaTCKLEJPag9TvLxDzYG3e2ZrK1X/uzUPVoAVjqxRWt6pb63H2Sy8k/Wgm06Z
WLRPl6TEbyYfMHwV2dtKM8O86yBP9NsA710Kv4N6Nucla73iK4JbWeOiZMtL5/5i
ThGcZy7IDXnt+KFzr5oX9ea5HrgS6WF9i0HZIoTW+jlgmClxczqn2qcdp9RNpE/z
ZFPA1OV2t4Qa1mECHm3kxm4gSjAr6+n9w5c5zSLIYLZuBdn4rK1H2WmVFdPFspEJ
1ZsWjceF95K4GrlSI3zV4IGZgUM9QShI/XHQFKo5xONiMrB9Z2Zu5HAMj5qk4iNN
P9tdNUpZ2sNbUHzWWprksqu6nV8wxEazlwYoD87PEEDtsf8QEXvnZzdOOakoovV/
wWfdNLCZ4QzApvrM/fPuTTlpdQUFj8cUANCDgcgr14MqMCiZuVlANQcDIu+J6mFD
aw3ouznGZyOmrkbJPUGShuji/GyP3FM/7zfG6EXcpFvhbGwHQJeMmK6xw9AUoE8b
XgRe7uysnOklxfH3eNYNA7yfAbKhu05/SDqytSzQkfEO/nz2D0lj8Hnz3S+BWQVZ
r98vja8ROLrfzH3oC2h9mZyao0zTGRkMus1WwDvSurAmKbOjj/SKsbDyNjggU6m0
8Huc7BNm4hKtcuhF7taayh3Vz/PSv9LfUK8A9HmgN2VSfMLIK29C86DTh30nTGXM
rlWKUI6072iBqx/YmiEQVY8peeuwmz9Vpj4aYc95AJOVvlwDVfVzbvJgqhzQ4Ntl
pXBaUvuFw2GusRqYFCpJsv28FergnNzz/vgYFTqZ6CxkIkXARW1YHzEjGB08jA6s
oEvdo+pFfMcXrv75MHAdixLe3u7o/XRgCztAat15fO7MGHFRuUpnVWukAq7LaiCS
kPILaT96+wgyFPfEuBYI0G9n6YEB3kS+T7ODowzWmZRSO3/V2gFkkb9091zfCqL5
a+aPphxBZbv/zM1A228ScSEgSa7uHEHPTXQCIz/zHrkvlSiS8yybO6FOCXhW6CQT
8twoTudy+x6eEHfvZrKSXdXja2+PlqMhz8D1Z1800LBDGsN/YcKRPsfNyIOZ6Eh4
OdhMPr+/VFszBTjb/0+ugkUnNF477tHWtS5dWvMa6JpzWSR3wadtm7NSw6pFsdms
fgCZd4XjfM8uPQk4pbM6f+kNpIKwNER0UUDHobpsNEO24AVi0DL11wmijYk/3C60
3PnDDvM5O57kVpFqn8TaLlPzmAxliQpMIiuN80+wiH3npHEUHRSqxaPKRVOvX/Lt
cajEHOCng/4+KfiZxlSJZRGrpoy/xyTEEJsx8mnNcmeZJcUb0OFcW0VxdcxaW7tS
DuKbDaiH0JgEPQaU0nEYohfuJMIw/IndEkSpwmOyQnHWuRgF1CfkFyYIsGETxusD
KgZr4vFJ7QcicHWMXbnXFHZMvoDiS5omXUP37vs+LZ1q7k3KVDtP5LoagEAo8NRK
wfdnHhlL75sXAPaN2KP2sNRcitAR+9nwNTyKEGRQDgzHw/PEW1yBG4BoUDfzTIao
TaeplCYPvUh6f+EjPtej7e0eXJCsMDMLWp4rrlCngCDI9QSHgHAauRjFUiDAogfy
qLp1dr9fadl8idwYSKmFoxI7pmOG4HFUM2vvtKgrfPWAhbpnTOOIcrTP6TANb+pH
vCgP1U3j+nTngTeSRvDbEOkK2oT+8dYTKsFUNqeD6R2dtkq84FQqv0kM5T0jTqrH
Bp3VYBugySD6M8YKt3Rl/8ZS70PVX4Rsh3mefUHrRwjirTzc77zMdnUpvWGq1Yu/
4axjDN27rO3HbPl+g77/KFZPzr+RpV2pibsmP6quSkypjaF83XO6OxnfgB8FabKN
SmprDyFjBbqFh+WOIbVfDppdBXZb/hqa+6AIUye97dtiDMj8fHHKiiegzcv05awU
BpfVaZ3GRRRtVE/fhSsvgzxOkpceZ+xCBAsmuCgni2f8Nf0tLANEXWxDdnJ4wELy
nH6D3iIadUDJO/fQxP8WV4AEkh/FjZojhX0MEwDB17dBWyNZOrkCRNBuEjj4I/LT
D7Z3GXDZZyUWSMO6d6fQZCsHt0XXPlw+U0zhpUh2gIbTz0/9AagONCn3gtDsVPAH
w0PwQGbW40OxoyPIMShdnviCgW5E2yAWPBZdZjbTwq24w7pubC5jTrWWGImxxtx2
1Y61Sl3K8DOaD38LKUcZlH/AsMKPqhF7fJ7zHAUGZTCi2fUB9XOm8VxnKxmbFkyA
DvQgnt+W328Memr2gRsvAoZV9SFvW3Et/P3KB8Xq/Q+jLmnKetucdesqryOnGO1U
sDAsCjmZO4YfYJrTjd/lAiovmQO7PT+ULBmaC4TenQJfITNqUKkw/Tc5WHpnOTVS
cpYecDDNiDFtWjh/m48HW67Z/8fmvf1XGlCttGxoHtcXNFok4/sVWH9ghU925uAo
3jPwSiwzXUIQxhZY1qioe5Y+x/P9+Z+k411eDARMF+8P7t2f7an3Sg00ZRFVjZqi
WScAhNKXM9nOnweXikN4SSQV7owRQSXB2m8GWxW86mQrQN5RDsKnmAsCYocTEow1
zN4mbFNWv9lq36VTtfWrLevXx8SEbAM963cL1tt6ucE/ch8Yb34UZQzSUe1SXVmX
ojt3CZwOW+jxW50yW8QO5uTT1WDvJOleRuYVTx4/urOBvb7Aq26IXNPgK7v0mgZm
Ep8LGPJQRiA3FzcqbDorf9DZBZC+DS5YkGUU3sj+iKA/WaD7kBwmPH+Vx8h6Yn2X
102zk005XzL5ualtj/7P5udFKkkvdW+WfecRGnOajfQSOrMfXf6x0x7ESuOkLGz8
HFWz+oTM0Mhv50uoeHY0wP9jhr0QnMQ4wSv+akTqfTMuxuJ1Uy976xuD+dLLZrBN
lSaxhS1VX544cPYYbjJBaqNRtJIRKMGH+fe5+bqErVN5k4l9Z3mTT9vcCwjkENQC
I/99npQMdBzTJfCiqLose7rUs9KroBBm7wOjvp+AYNv6dx+JG2VazAcPYUit3paD
dJW4DaHrwAeDUrTFhGi0hJ8MM4RWkvZGvNwKjnxYfXgmWPMM+da8cLAPicui5uJI
NvSLzIRCCwR5/2rDKusc+sRAz+3a2i2pjzgWI94ZhB56o4vGrbEJ4TS0YH6oxIwa
TeVi+9tNEXX68dYAf9Aouxtt4jkJ8qfTJImxhHD5XM2ahs02ADGW8T5RZnU/6/DB
ked5DMdc+Z58kOtYJ/PkdOcAyHgl4T/mAlOXaSeKSKLbznQZ64igroLXfO7rvVDT
X3zG93XEbLv3LzHd04v9iJVPe6kflczRKnS5KSZ3dO/qCaWaj0N9Ail4z8dbYFN8
iES71n8XYmFAUZ8/dnX9AlI6IMjCsMKsEOqzc21ab1aUeYopuECr6QIXWnKpRi/R
aLE+sEB4RnbtwcDRci5pTbtH5ApEDNNB5w1awmPPfjvLmFD8w4xqoCPp5wVjT6EG
dBT+D6K4eIKA0cBdZ8mJLu7DnXu61stqbp5NjVE3wx8dJUUpM2VhEwH7LWNuORiG
CT3dwgZTHNZERQUlibH/RXfuQjzuxJGvtAAn/oSzDyQGr19MZ/A4hzK4KYK6MEhE
9fMvkhW6ox3Bdb4uRDjbXBTH95Iiry8sObBRnLQ90uoVX4DfOVyvPRGjomRmJYWc
nk2cC29BahmgFOIBuAeyVHM8x6ogVWvCHvTD7ermwkQeQc457+/f0XPwbcY3fT1Y
Ig86FvYiHeE09nKun7sxq64r8ww4OCNxjaZ96bT/k+YdmKyPpnpdO8rzmSIeWWnV
REvx9+Mccs4Bgo+qWLz3Ra8kVH5l2IdLmTrx/wJEON+5bvHWMpSciQ1CrBwg86xE
zIibjGb2W0TALGGnVZuBajjwTF0sH/QKpdDuO5Kue94xhtthqr9wgMtMaFU3rZWv
hJvfyp9IODNXiI2yACP2rSKTkNgarzJ0FkjE5BeGM3hVqyHNA8OqZT6njDp1bjHE
IeOKudG3OS/sFtaoT+R4MsdCB2fsN/NbbyjEYjyLZvCFQ0Gg3/G8cHVsb/3jWq0i
XZL0s1g0l8pVL8q2ggwChKrxUBpRBYsAaPXe5vrctmr/ZncgDQaVzDfK7kK6SQ2o
6qYvsxvHEbhRwaHCLJozF0evTpR+rcQCoLXBZ3zWQPm6k/enaPoZU13Wy3ULJbEt
WWoNiS/irVQEUmGyODOmaG2N5dsIGc3A+6Ffu+62Q04/tRvOzao4vmx7dVCsj1lw
sZLJocKfbwMhfkp5jUmVoH3Tas+4eliEFJufk0dhNPuPoZtGlQU9BJP6nc+z2veo
5NSNJ4ZjtiqOuBDf9GNvixtxSsmyOp/EtDbPTSPNWUIfyV3rhpBudh2ik5YSbrSV
ZZ4OPcXwUJtRtE+smQ+w0KO9yrA4LHvR+o8MbiScIX1jHztuDwvrFSSHeVzW+UfU
JTEnrdTpQcvqGjPNmJitMVmqWqpG+jybr4EGszgTuo/1svyh9B3DRbAsqp6L5y03
dc2vuHT0GMDs7vnhfvrkhlOofpSR209Jzn0lXeuC3m4EfhLY53QIlRpSM983oK5b
c3SyRnpbf/FOCDqPfkM/Jf+yRcgegKdAs4yMGEQaGAEEBBJc7Rk/LLeK1d1rmIuK
Cb6ImD+4bLAipdSmtfLFCiK4kV/0MaNeuiPMBQ/JUvVjIZ15yDd7/gL9tbGIrO/A
VmdVqWN4IU4OTjOT3b1Jvvd5IzBpel+BxWSmDtHMRie5b5VwluDzONxZv01t0Gfd
9jsM2abxIek3nBBBVRLWNY85EsfIYXJat4JvpWZ+Fw9lBTmBDvyF3gUbSSBOXeZn
Uo0DsBgtzum7/A6E1qiDGlcAUkwh/v10e8SqrangKiaAz6LIQ8kWQ6l1bEH7JyB6
Jd9PxXxOac3kv18V2H0bbYY/mhjvrNHG2fm4ZPeKZ5lbegmtkSMalCvjnPbdAPSI
IFOglfpyveXXxayvNv7igbWb6ei7zx6ekgjY+yyrqekGX8Xz7S+kYvHKeq/+QwWK
h5uOx0+bMYSt0+xUYYyQ0IcB0cIdKjz++nsf5wG7RIdd7C8yV+V9FxgeScmzaaVW
CgzfiYy1UlSfTNt7Z/AOtgmbUakZRjoqPvvAEu1aFMltJvgZXs2+ienrsTuFnAHN
+KGLA0XmyKHUWdy1jncwMLE3FUVEMwxZK/Dlvm/uY2pgMblboJ/XHLxu+4mjAP1w
1AnID3cjWgOZnFDLRwLBAct2TZZ5pBeC5gHJbuxUrJqgLPVB847BWDDgPZDf2U8+
UKqGNMt09aYT37SfVg24eg+i0iZL73CxzeJhAiy+YJS0JZaJZ5NLIZeMEDn5MPY/
tDSdY3veGFv4X12WBv9w173PT7owRn/OABciUJlkktq5nIsnMEI4jy+KsY8qbv/u
O9Rt/lZ0If/0RX6JEan7MJRnKgGeYDDjDvMPQxgvmxHHTW5hTZopgQ7031HFK2U0
A4w/25IcX2eytK5dmMN8dz4FSnNxhuyesu4MUNtCDCQvt0nnOTxgxH3CWdIEm7/t
IJ9CG9OYFL/ULaTQ7pRA7NE6Mbl1LF7hqGrOiT5sbl6XShx8rBLmMT+2qlhFWWiW
LcL0Xu7lONzAZA9qid3Y6uQUai3Ao1ir4AW+Cmnbsd4fKzEhOKsi/TFs53qNgj4I
4I3ySJ/H+R/w+l3sTM/fmGgObrQhe/L67cPc3NlTGpCxBKmGqW6dzciGwbhKpfOJ
L7whZKH/TdlCy0wPkisoUWZcnb+XOhinrwHYeoFceU3cyZ4h6pi2Xdg7RpmMZsEB
LbabZwJB56WDPeL3dg77Fw38cnQpqag4mY0gHVfFM4yj60yxOV+xgV+1ER9rwkIj
4lT/KjG0kdS9tUftd0NIb2Q6p1jEN8ikOGK5Ei+5owSyigVCh8J5tz+QYFJmH1XH
sENZdwwqiHDUS9ph8w9D9p61wLgXgFppBPYx/YOjABqZjV8mqkXS/r6RWXq4ttzS
3PES6KgAkT7uoN3CQlPfG8fNqALIKtZLFLBe06PgUi6RvqJ07k5I/whq7YsudAzj
EQX1fpCEow2xi64kwajLU5i3e0fJnNEU394C/MdGvcPNmhLaGVQUbpotLbRK51SD
DIUQGUw75L5pqOPG+GIGLtdZzhU6HExVX+QIcT4p8VhnAo6MAl/XgmqBGZHQi7li
f6QTKzB/TtVyqd/luuBwf4fK2JUOZzdNYh38cBsGcpmxE6CLf03amn1PIr/3r3VE
degpVVTkIwztd9BrvmmIGwblozQ8sYpkEH9UyIXVSi5TauNjo38/GTYODIa0db1R
UNSjuHfTVar7smFzfgzQroPyUqdAYDEAZoaXc0BwvGuP6pWaiVNkxS0vDqklw5JN
IY8bTg8TgBI3nQvWzX3dByIHRLzAFtyJo3MgzTpRS5+JfSEOAdA6yoBWhL13/K7O
A6avQs31rW4S18lo/TXdMOXv0gfx4XffoWCjmpx9NmxcnLbJmKaFpC6IekSJJ0cj
ScHj1DKD5kpK9DoLE6iIsHvl4EfpymSz3FOeULGGjvpTyJdBNtHRoHN7ap56fziK
IuJtW6hgEexotNOtNPCBkidEOXbS61Hd71mhCpS8u4Ue86ndT4nrHm92dJJN29IT
HVfDoPuD1NHdpw1OMSvPDeqDia6nHIgoGKX2IoLWqlNEu2nirDpcYhv+XnyuNY/p
2q57ziLAS9sPEKI6StVKDVnXeshOhWgsaOf8IhhgDw7TSQaC+0QIMiu/3KytVCH/
VxOz2yU+Y8SSrPImdBjr2OPPwEwJeeUrGZdPz/ELYaQADMRtJcrdH/RnqNgIaGAN
QwHjUkRVg6et1IScTfctf/4OBcPWt/5Qf+yaVgpGcMYZNA4jEhk1qJltfXkL/PoA
GuCa7RU3wTx5CbY/eGRYa02YXf7TUIQ6O31H+LJXviGZpqunI1Yidro0w8lFfaCe
DPrUK+FsMK4w1BJ+DiurHvlOYl2NSLlMBD6GFu9NlfIQbDDpdO/K+W92TVSBRCMi
ihURPL30fdof3rAuRRrEwTT20QnuNIGIcr1OcDaUW86wqQyCd3d3B5VW/KeceyQA
G7qwW7jdNNlncl9Rt741sDQOvrJIzRyyHfKs3FKZGgFNczWwyGnuMCJe+QSfw+t1
6EL5RpLWASHzhI37GZI1NrAsANvBKmHwJu3rSsTQbFcZEVtddSdHBAOgTBiYFlCk
QlMHQzY24W23nd4uObIexgI0fZlCXJOCbADULsnsBccNnUaVXD2YSVTrD2sjUTzE
CCqkM+f/aQZmZE2/pfAQCbUiPXxQLCL/ps1DuBa0Y+bCV3XVKDYBPpF+nFfdNQQx
auN8tn1gxkDGX32vPjaZBHpQtHr6dxVmCHM3RH3L06PHMwY1cM8TQQWPQ3F3TmCE
kJvUeivdTis+3QSipQ6+EgUp5nENY1ZnkOMG0FJC4OC/gg7SNgvxTUdJRmtC5Uvy
u5Dy2usDY6hlE/8KkDWdVHpHCGo81M5VZC0HMgVW5TfOQDy/UwlfDJy6kmd2nuMA
K5401rlWzgBbivGsqhXMblC8mJd2rbu82svDFDekjShbnXjobbZZhCcoGOTdE44f
bFW/ED1Z5X1Y/kx4DHF6XWG45Y0k4ic6X31MmFwX5HIVaz3ZxKEbcx/CB9PfQUIm
nyYTbzO8dwyz0mNs83Noal/i2AVPwB/+jOkgumRtjqwUco/tZof+9E0dEzBaDLoI
IIvTntCzrb7kFIYnh/qDlp3qT1KkQu4DrQtcX7XUKdTtr7TOPRYHpgy5TlL03ysb
00YjX5HeUTQ1uZgv0Q8omqwhDG12avVAgo8ZspmNDxoxyn2lS1Q8k7kMEIvgCv00
xO6GVIyi0FIfZkjfAR/nKbUATYeV4oRwidJwpcIQQrna9PuEhyyAz2gFXq8mBrD/
BITryVum0IE/zDMPoBAT+1NYMal+/z7+uhRyNZYnwTfgNrrTzjcw9kABJJdFmPFX
EcIKGVfjk3BoaNph8f4Q1sNNkRflB/LsRinNBZ8gR9Sd3eFmG0qc9p3ewwj8hmSh
HE7qU2Cho0TVvYaEFN02Gg1HXlr+dGFGHVHmK+hCMDPvjru9W36+csRM3GYmGsgV
oPWD8bHqFKlAB+avLjUjyqmCsGZByjwHXPNG4ri88f/cbH3Ahsdjf+yeKuMDJ8iY
ZajxM2BfIwuU34C+VO5U5vI3xt9zbdU91JM4XtXAXEk8Na+MaxmXfGZlVGsl3ts0
oPAQ3NTfYwY/OE0kTEuDtoheEEsCOEtLeYSzpgALQZw9zNJDkVDSVthcgZ48smQ7
a6vpucs51aioBlMwrlWN9F16kOl+grReknE58XmpxHkJlFbjR5J9hLUWWDv7P/LD
DIIFne/D06niYXmqFncQHaBUdazWq+a6JjF8WIqRQkKDgSfkIOKtlaSQO4CSOi6Z
jsmNXgXxfYFp2ZRPsm8T0EG2BknKtQgxNYy3WMZhEeOQXyau4ZSjX0oFB0gUmzxJ
8HPVlb14ORXwDG3YrA6jY+ltmCXlQ1CmQU5ZaK1Ss/BsEGTqvzVXi9qqrjpNoyRY
JSiwIavjgZ4vGXJFp8/5dgbPgj9/GIcA0Bysp6HQ88q/7v7z2nId1o75NgYIZqCu
KEPKEILXTz09MbHiZTI5u7kXnArbDJb6pVCVt4lIglU56tZh1tOb9KaNUeEqefSS
pe0KnDO2HGgCDsEC4WM8mlwseqv8ksKS0GNgxLMiINVI+Dnpbitw0PLgJDEnYn6U
XW83FqXNj/vtoM7RVdk6cZOxxHHNqjH4MdHUtDunjeILhqMznxw+M/vsaIF9TL9b
BBErl4tnO/DcP5unPLmKlEMyZqY4w/L68RGbB/VrFfUaSJ9Yy/6rQ4AJYUAaPHbv
rURreHQDPMxk2ZZLAcXBboJgCUPV3INiknYGyTRivb5StzBN1dKyHH8LKAHJ4byW
dUMJ4GjkFzXfQz3vCGQh5pi8KMy8draEOQu6CtApVhznKDZLwO8GC/35Bt1R6DVq
FQyBseFg77eIQ/O0oTZhHIlKlFAXC8PyqqEY5/3m8Wcc67dxhdVz5zxiUntBtfR6
YaQab3HPZG+gf+3lh0uFCU1pPsw1QS6wg8cavVyc11S7Y05pUEKV5XCxBkuPjPzu
SA37/PtNyKuBGjs+RQanFzPud2tRjYH/UKdsu/XZcUeUsCB/42hoVaCQqzgJzwYT
SdHFLn9b4lsudjQHHoN04ZkOASJ5moo2siDS86fNSoZrLPaU6YkbQYLXP2EDRiH8
ypcPZulbgFRqYXJbblsSbHZYy/++jZrzn7ApUe/v79xBtsrWxd40REfassScAfQy
bgCT+ytoLIMT1M65EvXyotVrlOlmxsVDLs2TecH9CUnjoztbH7O/+CMuYIpjmzGv
dC1Yqz2t7eYajIz4j6QbhU/WSw5GFqHIDj0/lvjn3rD3W9nKf45wY2RVqi7Jhku2
jcqjnVvwBCz8u8HROQ5yFS5aOU6vWiQAmxzRWHMWTjOjsn2ICc6oWxMbDvb2P3Pa
QJzqeZ5mOXVTqA6Z+/uTTvfjAWrkGSzS5aiSzIPtUdxya2oHleBRIzzux+eqN4x6
ELmoMSXN7QdZfeRCT+z+XisVir2uQWyWVSQ1BD4v7w7PUBdn78JN+j4yJ+VOVLpk
I4CW5EAKBCg/WTfWLh47CNMgrikerIogzsuO9ySXhlHzJE3WbBCZbDuFE21e+RKc
lcomIq0cjjWZ5arplwDAlMYX14hxxZEqxRg6EBn8teKhM/hPTkG5+nF4DhWOgv5j
rTJt7KzKFHeIG7ERntatBJ0f0vpeObuE1xm1J37iUY8d4kBardLApfgX4a3q8EVn
nWZBmsccjclIpsqkPztUmxGhN2xw2/mp2fWX8medGJCp2kHolu+1cMXYC2+Z42mb
FEGVTViWxdxwW2WMG/wJ+1H1pI6BhSamKovBZPYe8grd5uffO7B9O42VI1EKQk2u
O2iJxdkJmmJeUSQ0ggi13l76wjWC6UiSkWP1RG9zNIP564KeP/g3cPMWoc0l4aQM
6c5YmmEB0sXj+qlBMBV3/TBoM+21lOVY9EY4r909abN9+5urEzMlVx4zuiPzxkaw
KwXwHGGnNJMTdjjbRR8grPKXvjCdZb1hWw3CJ5/a/PpUQcUhimtGDgS7w2Kx3xW4
Oyc4w64wAAg1Jic9v13KfB+7+j9c5kIRKwz4n0PuRE0xSXQXpy1EG+ryiWayaIdW
rJKCA5xE2B0NbFGVfcdgEL0+JF3RbATXqxBfhi3Yq+pCxD0pYlGI/d8FWpLCfMSw
RtQWzByOAG7SGwkRLUV1/BgBR9WRLgWS5SQiWjYfAet1QwXYghlBEuu0EEz6ygFu
eyhJLMfQ2DIFzfBsByTs+pzKEGK0wO7Gnbgg8pNc2FOu9NSRlErtCrKnEn/7hKGy
XaybITZgHj7Sgdadkj2FQ+SszfQ6EtelTQvMW+3MsYltc2LfQWzzL6Vf3Vv85miG
VaqoXjWbcZ04hxUKppWbGQOcUPoAUBqriBamf6Htkq5aTkx5cvZSep4BvW+Vo84Y
U/tdqSfi4q4I4QCvuhS80WMu2HerbuzlUR4zRtA/DGPbWJJYq/MSU2tvakg9jImN
p4P+EHgpaS7P700+rHwhRBuZf+qcjwfNnV1Yl3RgrP/dtqkXeilnC1T1FGKi11Wv
Iwu6BMCle8E+d8XopkqBHTSktD4ixo0VKLV4f8nBYxBeVnA+j3pN5i+noZ+12/bG
xT6TitGkex6KW/vrSMZBYUozxzsakml519KsY+va+xWKIzgX7J+5skYQGSyOF+cM
f18lgr+yhZIK6kyL/nvs6BU1qVHvYM0curIaCECnYCru7O6qQHV8k1ZCVdfU+267
qxV7XS3k0K3RqC8BXKLfmNFvepscs99KWll3Xpc+5vlWnzX/WRWqVfZeRBrQjY1o
kpHNCutmXBbDJkqo6Vmh1g2iw4fxr3X8sHGtkM2S/+xzAR9DEXOgoXSztxPCxUtR
rp0KAXIdY9m487GcvJp6MbsZkB/ZniG3chOJ0PK0Bo0hHRUu3aW4sR6Ji+VQc+WO
8JqHjmfwUDaVxHc6FCj5biduzcj/GUEvtEp5W7x2P/wen4L0PpsSDyGD1I/SAJS6
5GSwKbR7JdrTlEDnkW38fIz4L7c+yXc7oS9/38s0+wgIr5ZOnJ1p8PlAd/ZSVl1W
kS46FgsFwk5CcGT2a1Z6ANllI0QGNM6fgVL3QnoP0ShRRNNxzZ6g8m+h/dGcgSPf
U2NiEzF6QVUZPu2XLMyCjcbdoudCWkF90068sfafEn9ElJazXzBZWQdcBJjuvlwM
gJHNKi/QV4z0SGys2O/sOeyLz7H06PcGTl/Lv5y+iJ6JglNzKGAZ5wulx17xYeYJ
KoOT9xUHhBX6CVI8yM0Hah7dGVtG20NXsgjS8TXD7lUh2AICwcj6fTdEs9vTUrPu
QVeM2la5HboSRzcC1nOW9oBzOqhGi7xR+9h03Q3cebzAXH6UhKU80UCyRVlU6D/g
aRYa4vLYOW6UV/bSmMuIm/BDqP1GYR5pfgnu4M4QJVjyDDZpkVEZjptt7LqmHmE2
Lw751vVlk5cJ0hX6fOSQTKLWFlvVxb0hKe9/Cb0VtlQgq++6tKE86JRmSU3/BIcp
7t6ScVFNw/YGv7AeVzBWlNE+0lY6yX2IO3HtM2AOH9O1XE9dC85rc6/QmpsvQTkU
XDZ6lW9t6avkCPdbpH5LL5sVAUPQY/SRRFvFvebV9/QOzMK2wtOcyCPfCt0CLZ0X
V5vNVlicGtdMUgu1rr4MFoceaKhI8U4Nh+G/0Z9AOZXaAGy6OldUZViAfdmjzykZ
t4RBRvXaBuD1s6D4d/wGqxivm0F0kGjvQ7NT7aqVFeC55M03TXixXbHiVldVomnl
j3BpsFxAy0/KPwnH4Stknhrz2TrEb0TeR1Q97ceM+Tf+TeLqGq9gvsPl+cYo2kws
seYsaFJk8onxoi/ryx6VIUvfJDGoid+wCNUx78TiV3KlmVvaEbJhvcUUy8J4/EFO
0YUSh4mh6Gz/MToe6lRLIrVjqtgqpCqHiBivTZtFc64S0EWz2FvJwZbht6kEjr6R
CO6hBl3eAIptMrr34eAFWa+QrKVRK2xbn87rLOPJvzo5n7LiCT0w90awtbz3mHcl
eR5ZcNdqh6Z/pkX1YEZYPf08m+Xr6DWch6KIF7Yy4kx3oK+sEfnM5WWOpllAO0yi
96PvwnALX4C4saBLhS2akMCG1FrzvRlZpqbZ7GLTW39CGsDkRViud5XZk+aFlCK2
Ko8GOeBqunAyFGX6K6k9QtysQ1tOpVc2Hp932/PL/o9HIxgpgdPP68mWQvXl+7dX
CMGlF2kDU6JoHwoeq+11eghnzaZy/BPX7DXzc6+pQKPX5paWhl1RNhAZptsUk6SQ
v5f0MdOaMVRZUPDWzqYt+oITfVRf3mVWPZ76sK12Kit2ThJatUvuL3QmfRKJ92fK
MGh24Io82LNB6+qWc7Z/kQ5O4VpAD0l8xarFHuGUECFu1+HviPgo8gU2D6yuftz/
TTiN+6pBb6OmPsaqcnunGxwz80iiyyq9C6bKqS0zov9rw8MVYHYjjigHSsX5rsrb
7h7cCmYw4vvMDLArNpxRi2SimG+WH/p8zUnJ37eWaBF1+r601GdXsicr+655eV4Z
c583l09XhHVH/iQHm9wNvOEWhJpoynSO2ra2dipGyyQz7gPz2vcxphs1hLugQJuO
El86OjYVev+1Cilzq/jd7lYv4SbEAHz+jVD7NweuGUJvnE2HFDPV5lM70TZ/UtBU
5gE+hjsJusmKEAksJTpmWjZbZM9C5Z/ErurR7gSpvrLD7/ayVro2kfu3lmz+/i1L
lXwONOyPIX6O1YE61qnKf/G4azOb1vLbI2fovruoXIdgoGmn4wrkkBHqqzp1tLgJ
1BfHwlkVr8kLc7zcSJxikUe5/RUoP0VQVexwGYCKcp+gVfN8qgs70dlfgz1w/XAT
5LqhdgldZ4/guV3vDSr2Z3zsqi6ouMFhYrO+fmc/Oe+wjKGbB8+GcmQ+5ZsMDFlb
ifwMfm0O0cgpaSJBNjmgwzK1Mka0C4AgGImbUsGFBE4UckkgHl9zmxtqPrN3JHO1
MTGblReLo8R+P8kTl+clMDewdQFTCMw4iDV7CUzQTn/5Za6EZk/YL5tR/4B3o1rl
4wAzJ1svkHgZ0L0wijiUNSvkKkrfSwexn6A1mUIbZkZVhcYq6EfTtZCMBKO2e0Gy
tGOBV0tx0VFa8kCRDrQo/QnSEs9ib5Obee02z9NX4yOnjHPrkin5v06s5IJAID6Q
ApdEHJ/dhsw5y0RpSnzg8575/9SQ+on1px7KoeccZ+QzBZAJaV3wg3IMPeKbuLb6
7aiaeKoMrjXSSqjAPFm2bH0eef45UlsDwoAvwQjDACDeKJB3AQjz0g9N8HSkjHiO
Fc5SjvDAohy2gdJuxAT/Mfrheh/EfGRhJptf1sMMgNLtvbI3qbINmrNS9bjq6Jxm
Oj+de0H0OltwfwkO2sOqGOZAR0MrWSQ4rGDCcyGJ7pAo28FaRfx2f61AXqa5d5UY
WGU8lDXtsQ3m07qe4RVbG6+VR5sNZEm+tJxuvC+IsWSwHsgJk+6jsxHK68tZoF/u
OOy8TDGBypq20KkfqZtt+GuzpDaNoqvQxLBLk6ShX3aKyIbG9gQFsDAt51tX3yJc
hyOARrQqDMYXUDxBlAGUZFa9+Wz/mzCmDl5fB2zsn7swWlCxC/jxwFkKC748U27a
hsid9lBjqJirGe0kPMHRhFZjeH8lzis8dfgYWsAdap7r+ge+rryqX2iF+QPly4yN
+URP2jnFeblX/b9pz2wtXm2f1QPlroI+5WxLFriROVbMvpnnABdCpJDaZRe72H/A
ybza0quvfUl7/EwktD+zL6py2LUC4fu6GvK48cTMvllBYRWd5H4yTnrnvlw+TB5o
zJcm50mIFbbg25n6lKP71iGAIFS0dUrhm6IJj1yJ3Jcmnv6t/nqMZxfPnDypw0zw
qMTi2rkl8FEa3uBuu+D2eJ0lAL4foJjb4UCFSbt0XwO2aQgkMi7nUQTqZRFozu3z
iV1dtA9i9g+p8pOZBjwn6OiOS0OkiwB3s0hfwmL9RGBKOzF9agkmcFbp6nRCrWym
h8TjzSh9GOHybxRr/1u3QL/+20tp8kwrfrCGkmgau6whGU9ncpK3TYKmsFbapn6P
zniqfi/2mvK3lNGN8ABnyo29ECDJ4FxnknQ+HC5bCdWTpaanFZXpbnBPvarOTAFi
BIppYVtKyigMUEdo2YRfLQgz9UJ6wllzpVNx6FkXlnXiRbYGj9vU2CdUSwH0kj75
xe3eWOCDLJSIxnaCSzUe5puSsJNuBGFNTnA4qQaMHwe9JXsa0jC4ii2SCqWjPVUI
DlfNFtpjyV6pEoaec/SgLyX/3PMcFCqa4bonhTt1rh2kmv14YoTfmWD5997QV3TP
JS8C5l3MXGTGkl3Q8BusauZeIZ7kJymeb4QqQMsEeSSQJxexKMnA07OON8JLQpQV
F7U1BKGd5acknV9j6Mgio5i267wgv75PSzdHJY41VOIfmmvvS5RRy2cj/YdQJM5F
ziwBaZU1wSs3Gk5cGled1qYnh9m3iIRMtBqpfUbclb1OwnvHuZ96qEa8kP0Xycwu
EMouACGitZVaVkqWkClsdQXO9Z58qDJ9osGOJMn3Lgju4H35p9eR46rHicqloMjw
Mp5HzAPS21d7ZBusfv4xdaVrvB9qZlnhUofM7EoRv+nwHg9j8FwSnHWVONZe3ABn
HnH2tEgDp2cdHfuSVuFHRchC3eLTIUxK1vwk83M+/G9UGfstO6O8rz4BnMn31pK/
AdKfPz85+JZPe1fi9LghZVPldxTatBaV0PtiyMrvbZ518aj/n2m/NskN6ZSRX8a4
HTWFqtY3PaplpF6/qA3en+zzMP5m6jH6t0cDJp44WlAj2U/P96ZY2atKb94TrE9I
zT/HvaM0Qc1C3kB7bz3Zyyf7016Gh3S/+1xRZNYc3k5p2Pc8ZJnHSdC8/kBvrJPT
3qk7Ene8djydwhsTuCxl1iLJM30RSXWA/XghpCli9PlgSApmEk8r6wv9nVQuwPq/
XRdwciZPfq+GHf4aBrvP7p5Zt0zYZvC8DvtBaYnGBJli88CSUHoi/Ulf/Bn05PMQ
34bFmkkfIssejr2J0R5LB2DJoa+bBanVIyJSEU4b0oL3DmKH5Nhpzug1y1ltz27F
SzG6R0vDkHR+E+KFOnqxVH7S+uEa9XVusqULUYqHTbzZIIHnWETYDbvD3GflizB3
wrzpXy18/wf+lraP5RcVxvt8kMJVLr5903MGl/uu3gia14ivZQ+Zi4q6M3i8vA7q
tLX55/TGDbtFqkP71NVWPPGmMxN5hfpg85gbN35zWZPpNsTrzH0DPx4seIZqEDL3
wswROd0dQ2eFeTRV5bLTKjrqcn0CJfIvwAe3Ihg2S1tKFC/bb/TzbQEuJCZoF41m
FE8d6tcD6U69lef19a4tp2aKpJbMKL/zwtasCAcWzJOzhJkFU25FvJzU3mRFqY03
S9TbMfSS+cyl/ysCxECqpM5jA+tC0FFAOePQZ02ZByXGZhkEvdElRm1fgsA0GXt4
jaG6Vr7dX8pJZ6YguCERRlEB/CMtv97o3dExsvkduCbxgXSrZZ5IwQIB2b+FDva4
BzaCCcjqeriPWvizJTUixx4RstCBHn1ON4HNd9PZiqHjhuw6AE35aj0qkvsnKkFn
27xpU40qfNBZXhP+tFwZ539+NpRFaJIYfi90IiHMYOnAyl2DelH+2+MEN47YbiGL
HN1ZBYcBubcrztpRos1BkvNTselMoAy36CCRCoWUrAu2rvSQ/afEDIXug2wHYfaV
ePRzvFLZaSAS/oD5J31+39bDO4VK8DOb5I6ywXm7K9lSAtzqErwpv5BEkSjq3hJz
ZQf4F7kFE2XO2UKpu6ck51OKFTB/aaH5/kZU9MPcnCcGh2l/scqIg+PB+AS6HvXd
gqkgFOJ6jjdTEoZEJwymWakmC0stwAerirQN9Rk44lq+4iEMAurGAHCIad3nC0LL
722HCeglm1JXXZN6ANP12bT3Cf5kR7nej62LR5Mbpi2ZOz85Z7jNpFkn2CRg5euh
+JAPrpC+OKMzKUQUay4z5VujatlWE++zBFoIRrrQlOfOrXOhMq94L0yokxFtHBLs
Av524w6wNHCNy9Mrdc7HpNOL+3NfaqzVxr9PCqZDh7t347z955p4xB4WB3uqt3Vj
AMIbIfy0xH7cG/ciVdArDDcnfiteZ/kT8DdVNsD/Wqp5iVfp0QYrRtofOUgnflpr
ETuRAV+o/i/2WF1hDQgDiYZ14C2eN5KD1pNv3nXfa4AhcOeKpF0vYJAh5AC67Uws
C3WI6FnB47v1f7J0tP7CeaGA90TvASetB4C6UASfmbnzHjIrPgj9fxF9C8IU6LuE
D0S2+ttm+8TvbK6sZRvHxO82QPmFlK9+SAz56FjHaDLjZqNAAfZ0a+XD0SuRneGj
97ox2Wqp5CjG/ZcCi4/hy5fThQd3qnxezSFkOBSsoIwvZpEd93/ag8g1tP57/FCG
EzZoSpkYNVcaeuzZTmF8kZL4T5rprDAeKIYYiAF3sCTWGZ5MSeMV86FVLHFeBW+x
w6S4w8TJd4Jn9Gz6w/JD/2pwIrsTEU9bmGYO8UcsNke65I2/mrSolv1SOfYNmO6n
f0VLhHLeV1Lza2FaXLDyfzRs0e8/T1ml2tZodpnKgnQhOgCgnFLEBxQd+T+4Cgve
PRbaFZF/Dqpr6qPUbLlyfG+eUZ03VCwMxA1VHrlLy+yPIgVc5a60w6mdkLX1wbIq
+UA7q2uSexyUcD6ZlaMCipRewBTLyk/LnGced9Z8jLXPTN+oP0L8bgVRs/+FReZt
3ldVKxu8lzVfKLkgRCAZtDdU9yXePNAL/CxU3v/tnzgO9xkuOpGnyYCg4TzoQroy
JXxwSXr6BlRwDInmr4H48Y4kRJ6GKdqdt3hhtqFT7LxN72IHuUZWDt97LgFfYwgS
dicTUV+z/A83OnwCXuw6QHuNmP9y3DEdYAprCUC1jOhmH91ezGFJDmU1Qwe61LNK
LBeHZ4equyRJffNpNKqi/ojcUmAdLlyGH4T6FqV1r2nH1qRZyvthyeA9lhl8pe1H
QiG6QGBh6ejV1V49Pj8I0+UThlbHmR684isG6T1pty/WkbzbOGD3Ynm4NIxBYC25
Vf31u5X57pj4uf2eD9ICU4H0GrFxU9s8N44TDcMWGoLAdFAvw2IlvX6XtfXVZBCo
0I9DYEcA+z3/DytEuBst6+AiCMNLsithnnNs/sjd76mLJrWO8aeKJVcdcOSvsnNs
Kk+d/uyyJoKoODlXZLigM31Z5h0xxYj6BGUN42J3MKPZrbFrvp0ED8r5LjCfhjNT
oOq1hAnPKtikgjcZ/ht22r9qSGMB8qxLGh8XC2iTYsaqNx0NSeFwXxx3y1vSMYyf
mfOmsWxRTc6GURrI2f3i7zjPWu4AXKtRyprki1rye2Ph2BYfarncPNpgfDM6qpNM
bYphtRQoSVt1u9dB4N5cZ/EMTmI+VRDbzn+ZYlyK51Hvc2dHQq+HhhpiS1zHuPfl
elzDaafu2MRa2gOD0OeS8ZwWyTu6y62GbP9mKgFLweLyVJrcgfGCmHrbBbejF/a7
1tiMHk0cIYxVcEDoS8kv0YL5jr0IMI3ZzZHgA8MmrWUloB2Tfu6p0j5euEXioZkW
4GASyWzsHbP42Wmce3TPCcMT+bU1DiBOO33ms/jO8dfpNjHAaWM9h3WQnKzG2lbf
R2iiqBxefRTQ9Pgtu9U44iWNc4d3Td8T5XBIrOp5LIcfOvhYB1oWXCnX1YISKGkN
kVa/yZv7L2sqDptth13d3P2vqFOd0cvLmOVGS7NbKKwlQ/qOYUsayjImo/fLdbin
CErlE3bJ5BtYctcV/KRZ0I84Zo1JRBtLA9gP9kfwnB32m1k5HWnqBBcc7R4fXdfL
kYgCIm8ZJjZXn56sWek/rT7j65ciR2r2En0d156mZrFo+2HG+Wy7g1r2si8bEzhu
7aBckAJJh9DoXNXKz7xe/+xKn+iePW4BwQrmX68jmUFP8NL6rJEFo866lUPHpp4A
ZIBqPbCr3cGR26Kt7z8lEQ24d+QauGzT4K151sCHtwIMRvJvE7zSK56EOD+BKFVS
GzstP8S1sEKE7cbjJsPMaQLrddUmEsZ3mWYjDcvDgQXHOOaITpdmNMVNKOWCCqo5
qouZ2hXI2CIzG6IjsAABpobK3yp3IKPFkucc9zT9npEkDZxVNLJtNzub/ZEQDAYm
a3LqdON4n1TIjZCPyjTWh9VQlO+gizh9cZwZdP3Ar/gPkclcbLceTyArilkpKemt
3a8Ggp7L1zyALfvLVqQjSIAlxuv/pJS3xzuInRxFR4xmIhr7NZxPS2eL9JIuWcts
yfYE912B7TuilvSG7/zNhsAueEI+G4dom2kSsVItdth0UAa2GmJ/nrEYt1t7ttE1
keHgR0MTtqJI7zQassm+kIrRFh+PB/s3wTA9MMgT60fxoESEh+PTQ243gb6Yb/vF
FJ5AKs8YpaLjYwVpej27DVOghOUSwYuchEb/HBCB5I/y7osIQ1L+V3OBgZlt15z4
k5cc3zWsCsCBlk4Wv1Gp5niDpQXvOhBdDxsxLiBtF4aaI78tpJogfR432acahABm
tr/b1KpljUMVXyoLiv4La48WSfE1VaYTBnoY65QPPUET0Xanut6uMLV+8sFc+6ne
cCO5/IObMj/cs9XqBQeupKNFFBjWNCpOtubAWsmuW84YEjV1wglYkvNlU5oVSdXE
EGeWguaisbr5sgLpBBgOhzFKr+n21Vq8eWBgPStWMG6kk9mAobU/T6pjYz/ph3qH
AnsW+58HhpwWN/NE+pm/6aW/oldfsl7G5Ncp73MVD5cDn8qpY0RYMv/CwxE4fTw9
aH+2SY5m8umqoVmPTMdhDWzwv0jij7/qeIyQZoUkMOvcXeeHOvyx9ohz0xtq/SYc
o8KlC0P0alD6YiBzW3eweitoQ8ed8OtIqL5DEfJeZSckDFE0swUdq4LTEg6Z1Lsu
ddMQum5VHkbWQRIjeE7VHJleYyOfP2Q1g/cp0GXRqcKCS6wnnBL87GT6qrqYCb8c
5nBFiGMP7U6R2Ok6AfZva6/gXK6fknUhqj6qX0Sy3JotbYRHKaNDCD3tWs9mOIOr
ZTGaTCAWed/oIJw0tmAbXzm/REXfF2RN+1dJ6z77dmBuc718Qz9K2HitC+m7MnYg
dDtJZDA0llblZSPJXzsbQH5wsoe7hBNOOYTTNtabNCzwKaai1sCwqIaUK0gx2lFl
5g3yDxvJKssx+KWZMyebDR5jq62PY5gK+0SRYvhQhSWqoqWHjbFhc1uefD+cpc9U
fFlyi1xqsty7tUvm08khHvk76ZjTozdwInJSaXrjmZqR6IDSKjKUD1P260b+01Cn
s+6FhhiUIHUNBzI5ix7n/1JSEoLn/4xaRcVeVZ3u/ioIblzue5A6SmjsnwTG85Qf
s34pi+PbbKEil+n7u13HeeYp+snlcMCD0RLmn8qP5cQlbLaeizr6TpFGnOFGrnWf
6Q3dg5PGbv9WdYLRigtTZgU7A5L9siGzTCQ4XucBxvjKfHLAewmXBmlKhD0ILboN
+pH+RYrT4DNb69/qF1iN19QNa+B3v3BwVseLG95eFPbycNmnuMGQ+cW8MLELNcOs
DnB1fqKKm3ivBd8MBg4ZnDDLhjxi1UkjWVnozlESEkKmM034vzsYSOe+aXm1zbXa
2XoNUBbLdHbyA/AHVdWqYxezqaB75dnU/dpKnScAroyKDLu9+D2pl6JgNEklNMJW
0ARxOoOFLDJtK2rV0kejsJc3x/5WQyPNNJiBQ0OuDvJSZ7sdVfSnbpsfuG9rRjNl
VDK8zK63D+pHp6EhET040/3SlGdAopQyd897aubMeBgXnCuTJAPEFwtu/vp9zmXV
OPWj39OEdgpyGpb0dS6j1T6SDqdfKsj42KkylwAlYcgj1hYWbL2xvudShINVXcpi
Z5LPnQN4VB7UsdAhAlojLEnOJwue2CLjK5DdF8+0wzeXILgpgCkB7q2Ei5jqlDqT
pc1pDbIo7F5eKwPnDA8iK6izaIygpcD46jtfF2wzz4MzqXYaAzNkOGgx0AXFYYyB
ABxTJwwwbpLC0pvWafnrSJQxUZFTqauPexyHwIc/oLQfC4SQljb0Pr7Qg9uGPgqs
6mWqob3M4ZpK9DL/qHh2fkZC2S8/6psupSAXN3HnIgPRQ4UT7uMf/lewmtJWK1dk
1+1PJJisMfOpi0ts2ibyKi0+F5b63zSpKUPjG2SbrTSRxaGsAYxMYd1HR8MXfwTZ
1CUcDjZnUOwiS3co2l5X7q8fRTh+WyiX875KSHbm+6ujZqsExcc2dOnsWBNF3c0i
RW9w28mUwQbc4roGYkCh6YL51DTz/eV5EFSsbzKjpSegkg26PI1GYyTB+oSlCxhn
Ctu8xEOZKvNfNmj8kBhyF0ACfbQNhvs78wcm6LikvdMx8d6otIfjOCdqmHfTFAJ0
jqlg/gS2680FknZXU1SKzLaWSASAjSH+NWns28nbaMkDxnMqvafAFo/aIPBt5brR
cPWTr9up7kkcJdJ8JaR5PvV/so7YeXaGQ9LAHoWRgoRxONz64ze04a17Uy/KNtWR
gh49vkBOwxuD2cdM73hHEsjiMXBC6YMh3emCIoeaqlQi633r0pqsZDgD7T4Bz67C
AROsIbn0chtPtA0gqnrm5sC1FWMdOfCuK0dnRmAIUgubRUGEWUGIYlyQC0iopNra
32uI3ddh9erKcbgpx5FgvPAtfo36OCaDJrp56qamjQ4LgXLcSBwUSA7kFYOCnehH
95UaKUabPOTwBVf5yCBxFk+Jrzwq6z3bK7/oAlWkduyldpq10zGYdCmKhqYVQ2BX
/2hCxqqd60Rzr83Dar5HsRwJLikY2lGVWMXoeUtSY9g3GCCjhkrs7qYCp0lPTi0p
PtnP6mbEwI8wuYzb0470XzWh34gLFC70tapHP3eDP9fi9++l5EiHtB2KfENcyf0p
LygQ1AVbHnBk5rGExj0ixYENYx4bqV2DW1FapFw36ZhzfS94v5Q+uNWXmawwB6gZ
UxMqoySHLbh/STNh9wqVALyaBQ5/acADETQQqfOmPBlAQArmlgj2obFZzZ525Nn0
RzVdTdZXjTRl8t+58Da1asj9bwcrDTOKtugGKV9ooxVShBJiXUlKYbOglsEKLyP4
bM9ShB6brI04UjCcG1GXV2ULimCur4kpseAeKMLbGfBE3bSeONUExiYOLJv30pvN
2Lp2dhp+z53o542xHedX7Po1qx1lw6EQ9v/XChwBAKtqyU7OOuCSybGXJJkh+S0e
7yUa0PLV7beS1wpvHhH+wJrdwzSmlTTSJrrXqEVU3H0MbjUUGRc5HHiVxAa8/8Dv
K4xCVdQAPLMTY74SB/Esdpu6s3jT4AoEEiz4GoTp9cl175J5X7lVLJQlmmdIb413
grhJTNCjFUZ18YofKi7H0l23bdq3lf+oYc9sbQ+OLZE/ZEVjpx3oQ+Ew+8xftQZq
xTgxdUzdvvnNom/RbldqocoMHXh6IXgS+N5wRfHbGU5PcL6Sj3B3USJ4NfPn83nC
SbdVkXk5cokRNMuoD8XRHy1b27r2Hpq2q8N2JWjHhAD7KwSZfS9YQuDXnWNh85zK
iPbTr/FInsMyeCdTHq19qxtgeSHKs5kAbQPhN9R72DQK1KV/cF+pIv60SgiGBais
zj4iAn4fQLVJRZOzraIm3vXJV8Aq2PMD24XvYC36mODdy0Snov6O5if8s80b+v33
3cF5GvUjcEzNZnhM0U4ZBzGLXykLnUTBiEnaNXUUswAfasNjOVG45W3Jffm/glNJ
KQpHW4Amr/No3U3dixnqCDEO1XTrQ8ZZ8EajEkuq85kFJ3J21lflcm/pLjKuhcBv
h2FW5BROrXFWiNdn7OragvPMqt0YI9RS/JTMfxRDuh8k9lDcXVuY3B4ExN8Nyui4
zbV4MZIvF3wuqxocZjHuJIjUgjHZDg8oWwPPKIX7CzKDGjz1RR3w2JF06fxWkSME
MHGW2+fAoRfazxHHibhCRzs74KKIYRkktsCbwJ7SSorS0LPOVcCRbC/tNUKhBew5
tTlIRaa3wjuPZhP0eFXRqbu5cmkHytnc64f7kgc/cppxpe8nSE81ahHj2QuYJb7V
xVdcuQrgyfeKjCdxRGb+80GpbmpDoIajSCTfaEOCbIgwIBjqwm8k5j33WQaQgFAw
gP9fAvkYdpbi8CpAtoNcKJTWDIJr0dTYrN9aNlYJBcCEs5TXBAx8RpbKnJ9q+n/X
5JJnXqazbSy8ZHH2/VpQ2RiKAOPxwQ5Sr0ChPDFFOjGZU8HNq3P04usT8npqS2cG
MQj8IfHuHTvbhLPXKrFU73TJgAivdFyRKUuRg2vI7bxNdA44inHIQ8B+Sfxriv+o
NFt3R3knvWLwM1C3USNvB+ttI1eUinGdzGJqH8WgDvrD2alYRxnqXprrhDgQbOE8
t5JkPRE0yb/v90P0R3jSii0NmCBy36U0CFnflle82XgKc+oiwBAuVk8C4uEo+Rrv
1U+DUFF2jugb+1SI4KzxfrrQc2GHkMWxLDQpRlIe0J145awlERNcQK/YhLQotPpg
f5q4gcbnqRDBMnL863fBxbb0XkNONruJUNnhGJFjB6eyaMYnQRXO2EwQdoSoPz9x
PrEd5XbEe8Yb6RotGBaLSF3Dtp3qfmI/vhhmhI/Tjb2OWmHDHWoA47g48utPEHIb
nXHMAArQSJd4Zz1DgO9a9/PqZqLywP6e20RuNoINUsW3ALmxU9fenZ1fIpvWpwrl
6Wt70HxSQhkdMUDZiwTl3NKc71T5valil3sMnneV+SpZxXDF+57rtS+mtbAIVYvq
rbgusj5eDsQYZM1WYn5zKcVW/g6uM2wFkUCDIjv+wjcfyhd1XHE1UA/i7Rtf5SQM
2GdEldHdY++ztzdYBzMDJcwJMgBIcCZ5X7bAHRKCMd6JF2NsDOKe1lnD2v3Jqiic
SPzDRV/ONCkCmC4n6D1bk28KbFbN3VP7fwoB/J7HqrdqWF8+x8+EiJFy3zy2CIu+
b+pTY1rsAskzKzKUl8kIVZ5XFaJ09lpu05XYR6Orc0xUJ/KNEMqpgE8fPVeSN2KA
maLse+3G6kDonlwriMrEx3POf5Wr8GRfnjaoOhksyGQhH2dU/PcTFUcvnYZbKLzC
FVdJEjZ2frfigMcBHYLKsDt/9PD+67M5PqXSVxOCPw5tIwfQIiq/uGv2t4WCL4tC
y6DYRjYjhmDQGvH3PawqYqmTB/BepmLQwNJ0khOo/AVylbrQ/bHyO8MnkL9sHr6S
bG8FyuA4w7CuDdbzn4hU1VB3nahOupw8tAECFm3bCBgfKSrfAbHzl/5xumtUMYbH
l+RN0pUPvbVJfC590gYP5pT6rCtyua57kkLyrmsn826QkfCpjoHz5LMhRXYf4TG8
2WUOnI9e5NocUxtbwGAlYvAPLGDornAnrx0+do7pSxJ9PoVel2USfQE26uivAHjl
qFybuncw7rMMLWkrBxwfAEzrwqVynpP1uwrCcHlVLtkXtMgFSG9DBd+sH0oovjjU
YSU7v/Hhk5IwjKx7+LQllcWn63FN1TX1LId5EuLTItpU8P94qqYoCs7JIfp70faW
O4zwsn0C/f7iBEY/5v+kvBmRJg2VBHn0h9507nGeEclpfUYJUWEdnRTXfSQCgREZ
bYW5aJNuR3OFORO2Eym+80oYZ8QQ7JmpELfR3zQ2IqRidAYl0mzD/AEw5vNGm8Dr
ATsOZdLGrbhnOE5fpF6W6xaCrD9JOzpdhUKZEWumQIvPrTMWOR6suMkoiiMhG4RP
UYBuuuxMV0PCphInjEC7EgW+l7ybxj5aVrgNK4OOucIJZoclLwLbRH3Z9yuvZCdT
BbFFynIC3C65G9H5iBxoAjA3aAKEk7Ijmpu8XWbxY0chmc+4i28hvJXA4oEO0/Tp
TVL6QekKGZFsLfze0EHmwoyNgoFhf2x5J0CRvLR+gIqYb0DzSKZs/6Ta96Exmq6d
LD4uwYvSIIhuJOS8wsyANc+33LasLLuXLUkOYRXCUMsu4zws4tJZfS5i+eQMw1PA
+exgZjCboDLpEcW6Q6hc08EBBaEhXw48r5sR/SgsacL9K/0oow/gIBuwAPBURpVc
EfcwPCKwcyIZbcjQBtiFAJDbp0quzNpE71eWbPv4D/r9nNTrQ8R5IUhDxcW6OQ1u
PWo6TAIV9tEBSLl/QZm5a1P4yhGY7cCqsAGyQ9W25VPFnw6NYfq9GIm045vBFgDE
RfChZfpBaSiFzINIYQukqbZiQ4kwwhicHR533/JNYG9buTYtPgg+T7KdKavPl07F
hENhR1vvpeMR6ZJX2jdIcqn3GfhoTWHicYWErspfPUAB56L8dNFS2pC4qfY+UxTl
2q6ldNDLUVzk6pXWfKoUB1RKQC1A6RIu4vImBVZrffBE8OIbnl+XlHYlu1Xuqfoh
LaBOOlYF8dVyWHsDrnqsu/gzYyk5FOSF8U8v26fZT+2Yicc9Mel43OgjCy4VW1ne
n4e5qTMc7FUdAZHrHcCeFc6qyhNeOnfv4bE9GJsSc4nN0TPXKJjiohOz9mU3qc/X
YKJppUF8FO6i4TALy/b9h676d4hrz2hwRu9ap3GmWH3Kir2E1tIAnNNRUmfyuMaM
tIAcW4IJfu3k4SpsRG7/UYdWZcWRNHU7QL3bzERL1LxV5d+e+NXBpLcQrL8VinOP
sslQMVQvGZePA8q42WGfPErEDW01W51J541mQsYxaiiBUdSXOpxogfPtT0SGqH62
ikm8VSFDxAwHPer7+WRDekX8hunBemM2qI/0asS88bclUXqvasln3mWsdiaDzOk4
lLjqVQthrg3WY0+u/LfP3vCioSbw/xvu39pgSQ5Btt69xM944MCu2c86RSa6ez+n
yjJxtbC0AIbTj0LhsBwYk+6qSEiyMbNkmLs9Rdoot5Nq0XKREQL5QyBjd5CN6V0v
6ZvwuBg9iNOQQcPCiqxXAczu7NvELvWQqPdXtEcpQV23kxCMR+L70JRWURSWmW+D
9QIHWAuniPAuzAYlMrnFrG2cFWE3LmQabwUtPfTlMoivKxwzBL4hsGYP4g+e6jJK
7SN2fdeAK9xeZPH61k5DwM73V7J9HSAQaEcrsj/rgcy5WrlSU1spTbWt/pWfvRQR
Hf4+KlOhZrziOomVa7n9uCN/2/SmYGvXBnaLNqBx4VghDMZI9MMgo/XpAIeSuhik
Sfuzc4lb/0WDoXGfbM7WJxBK4iWr8aPigcPBvwPb7KOyyNIJx3nxS7sZlq0vM4On
xwOhZzVvVkg+5m7j5JjNUE0uB4I5OuGyLvmZRaIhEFI0Ej3cYeT/k76ILg19q2nI
dCgvDakFWkTlucrUZYryKTuTzyjklqEvwDMUbWZO19xh5GvL4kbWTk+JKc70ZSaH
EXEJFIEKtbPenO982Guz+WX+UCXQtWzeWNkaQDnvmtn+kLpp68Sczng5a73+ng/q
+qkpwgabrHTaInwcv9kAFAuaAi5soS1KY1Szuiu89WU+EM/Uc6wbTzRFCEQjjTrx
s6p5IXKjqZPK3ntNadyaiSUhr3H9A6ZrHNiQ6XBV6c66Pgoh/zPRpujiVgY7xCky
IQWfPVFetSMteqHgT/ZcMKq45XFsUL9U6D80Dguy/1TEpm6nidVao+5UWN4pMOof
VrMypQ0Mmkg9Yor/Lz5MrjtcC0PIozflowub4ZowLjr6hk+w2/bzNuA8jtsff0mF
Vr9A60hz9x7aN1cqNVa1tr34PYU9iqp7Rzwd2XpzW/5ZZqKD5qLbUDOWI+MD2swa
4g8qZnu38uZtDLawDkqFwN+AjlBt/sCyNmm5RoGG/ZiUsotUvOYj3/FhOz5fD+RL
Cp9jIjyRzDkLofW+iddx8Q57gRXYfRDKwjDhJAkME5o3pPCBm0OkszISLHsffrop
KnSyTbCJ3g+goxXzkFf/7vqNiOcVBR7IgynAAInVihQxcK5mYAXe5bg6O1U8ZVG8
mYTx8yjlDi7y/yBsl4cztQ1+waGLaeUxaHKw/qC+eduhQ+VeRchaf6flJmubvqLD
HuM9tdIfe2XvEu9ZGw8MwVNyFHHYkJ96NbJDbMFPLuvSVo6DNYrI4LYEYQdzHalN
VNWey/5hhzcxSIYgeg30sfkP/odlBktMSYSF5zuYWDCgQL8Uu2CAXzPKhDDCN+X5
5ht2F6hUm8OwBq1r10bGUNBxLpbZIgcAnLJlcs+muv5nYX4sz8J6mdS9M3JHU/GM
L5gQ4y8ppfCDBZU9RLSpLmZclje1wO7v8SS1tuMKudoM8RVlfAG+xQ0VjKK36Z7K
I0dL/H2Y6Sy3ahtvwd03r0h/aFl6hAgGJgVR0QZCLyCxT/ZlNfvfk1UJr1HZ+E7E
+UVyX0JAi7Sey+PiOzy2h1FlGV3NHagIWCxUuKnsvpk7iWoN2JFDodRf0kwCP4uL
cwRqzcz9Ptq8WOK/Sz/JlzFl/5iSh0Q2UbeO3+2O6DXGANB4TMF895sONJQS+3cX
VFF4orK5R4CyeVhZPRAmLKulxWS5EKJObeLqfnf+I0EGQzjKT/lQ8cZu6QKzT3xr
gODeDIniMrD4Vt7crnOvMsofvnunpLKPOfgDGVkEAhDeNUJCy62oMOBGU6kO/n9t
Ix2f2nOBW2zqvK6ZnfaKMJHGHBp4rECLMa6pKqRwZCdSECis4VZWjI33XvPoF2Cf
j71+xW0MRD5dVc7piHpNJhM+yzZtjV34mepxfqPy6ATgLJ3IzZt9nSgKk9LAuiTS
k1qnlKTzfLGPjWZN8Ys2on6l59KoTL2INGpdhH1PlMVw4ZG2dk/7A4zAQqBRk7Lh
wE1ZZu2hl6/v9PcPSR6SLYlpS3qQcKbjK47TbV2sTl3V2GAWot2ps2n6EsvLYGhL
nMf1yxWLg0vGK85AIqNrAMN/wHlehUzKIt78RCBqpiCFJNybqQfttPUogXcdREOS
KJmk74s/+Z6nd9MtydeEazNjjNTTTUPNvB54wvdNb1B9zeMalqIZv2JgIVkRCZpH
sDrdcaPN1HZdZTVvhhrnjZfUBTg2wRHc6JDXnwoK+J9XMSpWspzmXiqakINkO4XC
1floumB0GA/4bz15fetscWlrp1Qbygkz9wruJWOj9dds293jeFuYDKNjk6bxpULU
X07LHCcJd8wWBNfc3MZH9rIc4uq4/uiKgxLa3IGHAvMMDGq6gTIGuGnO9O+qpnYU
rF6983cOEoSN3/8DD+3IW9wSJR9h4s6cu850fxUgdYJ6xw6ObTrYKhHx7b1mn8go
wwZdBoG4H6KrZL/qY20qMGNmoN16lW5sD7SU7QHwuqN8kurqoJ5ogCRYV27mrjwO
56Um7IYO3QQ9lNYbK2YoyayRVAB3bfdrJnoTv03pJLVxRlH3o+WBlq7YmFqxHJO9
UscUzI2H4EYO+u8JFsYHGpPn35kJFSKbaaPXmhOLO9hsePB80NhGWormoLxe29HT
3J93Rgn1lfyT8nK0h/GzIcHFuVghHEnrppqnFZHqqIlTcLpU8So6wofKXslZLmTx
elEEpsDgFyGB0Bm5Nu7p5LtHXEQwv83hTDRXoW7KQMisMvkdR1vKSfHqIX+y+L8E
T7FKs17tHRzLgMDZaOW1ZQPMzmVidtRZaJp2BoX2tMakJUoXHn3oszKz56Il4RZX
MyLPwJQAQRkhKNa8XZ5+toyfWC6j/4+EJ3B0G+TU1fRZEm+LWe/tw1B7CLni//tS
ePkVdO8rSljspQUAL03TKmagfZqJQxnlbyyyh3q4Amyfwf72/2kU/NR4RFuMPtCQ
JttRD/Gq8m7tSUo6tmqGRYOxSxqlKGmZ02MBDK4Da+Jtpy7GkcgEYmv6WKXOWyp5
wt4QDg9OWYmE6/Kkak8b6MM/iaI5DwNDH0t3he6AvuUunV7TBxxM7TsWqOXZZS99
Jfm2Ihito0lCovsVvdkg2ZTXT5XicHIgOO7kwMv4R+psASy18oloBfOeCsbJfl6F
6CsJu5OJzZC9iPK7RJ47qvby6CVDpKRKhB2zFDCZB6N468vG/9x224s0Vo3L7Jm7
ch+ltVvRyn9iR+N/aR+NfhomUPd7RxzMRp+wykImAYaEVS+mzlt4Hjz5k2pI7hQQ
H8f7802kNePQiNhYpEHkW+oxrhVJupbbZK0kwXA7yNTbDb1wjQDHo4a9vBFUC5Vj
lOaqXD9I+DpJ78l4WnDJn/Tx9XI6OB9RCRVt8Jgh+1rf9AY5Xg1lR4S/IbiNlsij
v9beHsPenl7jMOQkZv8XbcMPUX+d3MQvCwZ1+x8oFbYg6OI4pi+JgocPhIHeRgUm
hDBOq3ynwCS8p1D2hj1v6klwPfdHMFyxEC7qe5+AMJzVwHN1UQb93iZ066+9glvp
r51wzMnPlve6Oxl67Y/OKDjlWCqkNV8Uy0tyW3/0lEleDKNcAkkkzvWvyOvGjZVp
aWuhkCp3Fvr0RGkZalmiHcKJc0HMyBUiZx/jsCzmqVS/tqyTxLZZW4G9OoGN77Kb
gO9uLgGDhyULqyfpA4FIeI30RtjRq2KVdMM7fDsnlhSgTgwSgxSU8M2pv+yCQIsG
sNc+W+tuJxNOVyYLj/+Cb08CJVxBlaXh3XomSUT1BAOsMwcoa8IowpgP3/iTk99w
dwa4moOWkWuplhAhllcBUzmiV/1ROMkvQnwgz29AOZoCqU1NveAYEaa7KZbNKzyU
fU6Kw06p+0+GDg1mus4uNUDk+OGDvA+iV6wLfa+LYJoDWW+caHQrtDRMQz6xBl80
zAjr/h5WwH+LYCw5obBwgkqrC/n8eA/fDyEeupuPoqAY9bzQMFupfPlyW0pkGHkZ
yx7adQKvlATUmaeaFGYhS/zjdgQiqZDlRvaNletY3y7cZjaS+Gn0ZrvGEbnXFkKM
umIZ0XtL5uQAekerGbz43wXA3SXyWucQ4mBX4dPxj0Ozdk/r9LVjvd/J2zr2A1n+
6Dd5lEm/t3qd2oFMq60MCp5HeqyqLHcoTb7IX1RMCZELrE5PJ+mEdpinyzkPtG8Z
8OTyWaBUm6+NXNybIixfvscatXR/VTwnMXL6bu9WkiMdXV8DYVov42LIwdolNeQa
1wdAvO1mObANZVjNLLEN7di9tXc6f8LnWonPWQmhwGS7POXG3+ir5HK2klGa67iK
27EnX940pP8limd2hkotSljHYWW8yc2nXMfOoHwn7o7Vf4bw0N4ClQRNFeTKEg4j
MZF1h7FqocYYiIsozL+ZoeetWCHqV1Z1ZTWb6120PsNOlZEHoHa5yJpGuINl5wTd
IYx5DvaNbtqQvqIW9AMj7WNpKv6FjIx+4uHYSA7GIePjmtDNkzc9mv1lzZEmNV3n
t2j41K6LGpkFJgD+6S+8Uv2k3C8XkD5wT+06uz2ru4rqKcfty+RDEap4yGbmsXLn
TvIF5ZeQUUe8RVeMQPuChr4KBq+Ajm1VlPv2IJBVxHmLzB0bivPL4yv+lBaj4PJ0
oqYSwXChLyYGCTL9y3CzFG8Wdb+qHO+rcp2NHqK6luk8TkoCq0EwDLgY4zfhKCzp
07XV8rA/ZDJBw4trGHeuz38AOGfjK+3tWjoA2z2+e0LqcgWvL7izmB3jUmFU3NeJ
1t2PGB7EbodDDWUGAs+rmF18xYUYHrkLMqEFKc/iO49K4hbUTrI4lCiDHd15OD9K
U4o/ufPvTJFODTq1hRN8kaLfbjaYJsE+2fcgkb7zAvQW8iKlRL2H1UfhzEbADVpI
HHhbnDSbVJYOqfeLd5QSCSd4l8APA6OTipm1e3WjpmJaWk9mHytbV0QEe+BK0fdj
2ei4cRs03zDNhACddwSNTAz3tLRqAylZnSaP/aIVrzPCalT3HxG7PCW7DX29NVzD
kSX3S2HkFF1LgKcTPU9Dj1D9T3054VmsqaI/AJl8mM3RPduXK6ss8QNsKfVCn/R4
DAUMIcZu5V3QCNU49bYOqmzT76Whkklfqy5m4qzR30ijlWqvO5k7ryM1JTA/Zdcb
er5mMNUvbSE+Owr/qA6QzeB1zKkCm1cedux4B0SSdT/OJvsfo7EfCHWaiwm9NloJ
uFDd/QJ5kNQ06bywk3Kz5qZj7ecehqX8G459sRt8GO5RGN379WpUy6zVYixzwu7p
PC0d+jv6XNFHjIU/Z3UO2QpcqBLt1Hu5+kZg5ENJn3ymSczt8DeCq6p2lCBNOuQe
1n5InevtKKW41CmiiR4UWkoc4N6Rf4NEIffcKWdhH14xUDb+2mzSk0/vJDJCE2ad
UmA4e22ho5zTDn5Muglj8yTW0CVmicu0iUOzCQHcc3+ek1XVTYgM5pJdb3GH4Gyc
wwZ1T7BxneDyQ16n4wDjX8YZqrUisXrB84qoW6xi3c7A/K4+CK+YE3DCRE7YdpyM
JbE7cm23XM1H/J1ymlCiisRLMqWy+/4AQ6kZf8syTh/gKRJd24kU1laEtctd2Zs7
QhH8Z8cF/lDuWr0tctt+mYL0qah7Qna0Fs2BWESujRf15tGC4x5aZpGARgupzHzl
cD5+QLy/pXFq/fmjYkGxVEa2edBNQTQOlK6CnJ3wOpDyyArD0xkeP8iyHiNjRG8Y
i/HmHGwHjh9r0OhFIJ/yFb8LMnew4WLOYw+PlzyDpsHRAP219581EXwMSHPvDX+G
ia7mxMO5RXVyDQLCiAPiFeIuGHKd1R+j+OSqWdIQmPTP0aNI0V9fjUiE0vJyRKOq
XGmGUMoxBiDXOIdIQJVF66IAbmCB2xCs1cO06UWO3dNESXDvL8synX7zyvNiZ+O9
2Uy27Hjr7yQlU89fvAL5/6sHVj0KEh7KGX6U2DIBFpVHBUWJZKKH91MYFnyQbTbL
vHb3engDF9vE9k89fONoHTK2I1r/RXQ6AaxLdFoQDlCwnkSjCgdnSq7eBFMckz9v
6ZDcVf/p0c2y3pE9K+3CWa2aCzKM30HFC1dvIchvcqrohcwC89/qpj2yf+1WAa6m
bqZE0i4rU7Ks52INIPBOP7x1HGV2Lbz8RNS0Vcvj9dv3+KTPJ66fQ0jjZ+SksG7b
VeMLJ5fqVVgk253yuuamVp9kgMI5e3D5xlVgawS+bzkldkPL2nA5hg+5WUHELKit
4pq1EVDDwNsAaZ2Z/nQ1I35HKyrUZ03qqUrbLxne6SXfJVWEqjOJ5TUs3yBbia6j
JkwhBpL+gWsTmMx8avX9hIkY6bEQNeFdAyZjK4Qz/WncQesARYpKlcnkSENTUza0
SGJAkeQ8JaU1IO71rqUD4XPzv6UqNUx5hQE/yZI3zExQrMg/ZJsp6Sh9rMgj//vV
+CWV8WGS21R7jZI2/pps6rqwlH4lYeIZqtX65JfXxW6MFAnf6UdC/KRFUNYToSOR
J80cptmLubCpJAKZAv/jTtZI2GPmPoUQ+QpFBu8ewylA0QHrcZ7xVAbwNlpjdFOG
9uqWKdZLClVKsmiTHQ1F5BjVy9pj/4OFeU6wY0W1mfRnrv7xLA+69W4cViHbtClJ
wG5Hi0mfnZY7Rmh1QqPBW968QmaQuy33qf3SP/A7ygylVruHZ6eK5rfnrUSxqN+1
QKHF/j9RKgBoTIDutTxHqmo0ejoU/Izs2BG+OQftN5L8MU+9SHynsKGmyLj1pRms
jMs7kExNYL5+G25JKrOYkRYzSOsVA5pii2rHYpa3OyIT6pNbty9IPtWhT1eFfly1
/BAoybvK/31OCTVvPQMiNAsoH1W68Tdsrf+7OMYeaFwn21+9XpECl5KXkcFc50Pw
o6RGTWGDHLBdgX3QBoGiUaNgg+atb4YhROLgRJ6mi+cuU2b5PrD1CsNu86lRE/JT
6ptJJ/yrt+0OqO3RDFTop1IXORIjPni4McoV9qMf0CS1cXx0BOI1Pq4TGO7R4Oz5
heyIhEPw7bVNQhMRZDeB+fZXdM+bW/JtGJWqSEYXgl+YHJozXMP9JXhDCpyuKNsi
yaK55psoFq60fmcWlLlGSKRcYQRZniadRNjxZQismJ9CQn4aAsDT6Pjb8TFGjuXm
TT/Pt6yICFf1YA9/01jeydDs4imwswd9aK0CgBKrt7UxJd8+JDM7RKs/869/hV4q
zSqNWcpdrfLk/KRJxivqOUr4T+j2M5OG9b/xNmSIb/aF4BBF9EYWYamOVmjhDa6C
tzVqym+gZ05FjdgfLB+EhKuHhvQjDBsfL/Dorw7UmN7/w1eQbJFxehsLqEDf/UTL
dF/dnLqaj8kkqh2G/pFQK5y8IRVTNGaJPSCjNzuwZDYftWtNhXk8z6KX5I1TNqQO
jXJVWCamdNg1QT0dp6/P5RuQxsF2qIoAqxQ3dhdMlESJAHzwgHS6hUNVcx1XxL4X
UHywE1bN/RNGDSpC6daR8kQUpzUEYIOwSjmO+jcCz2C9T2T6HUchOHofZQI4BlWn
3vJsqZoL64FbzZxBQKcmbtcsD4VfIPtcTs2pGsyLg+mXh/OX8GNm4eti2LZd9LsV
Ho56liJ7CXkOvYauWTgxoVFOIj4I6ceOyUzHw5sq0M5k24AmvdkBWGmdxchvf64d
Nx2QwlW5qA3yLbB6uMuv9DnyWGlkL1mLRliNx8BU5i0oJjyCV67v938ZePHg7Kgj
NL2hbTXUdhAx1nfbFetu41Oy3IcmVKhKPlXOizvGTHao8LyNXHpppLYAU0Gniaun
YlgMtnVohVarwREXWEMwvysba1OPPGYjLCamm6HcXnipkH2Skg8TGiKIS/KIjuLy
r2lxgzT+QFzo2zVC+zE/QiYHKAFGYSSvflsWv7Rtpres5Va21Q6HBYla7iWuFrjh
8A3MASBsaiCAajUIPm03URTd9W2TunJbKOcJ9BbUAm5vhF+vDersZOvE8KFbbMf6
Ufu3hD/vaHisKkMm1tFI7l0G9fmwxBOeEFlMEoE7DEm61LCrW3lh9o4oe0TxT2Mr
EtqQrmqpO9mBtJalSpdVmmZST1WTGhX+jdyGNXxIMnDzqmF13w9yMyManikxsvwR
2p6BOBqb+EsYlVH3VkHSyRvrFq69SoNc7qFgPdlpL53JnM+xr/Cdt9wvZQQyB8X4
UjmFFnC47sj+O8S1eMh1o955OKYlQ6eO/NVrjcgdRvX/GMqE7V0eamX+3/JHxbwz
D6wMv9/mu+F6GMkjTph2FFXGI4MkLT0PHsXRO6KShXglU34AzMEAfGyucEwEtNko
7WQyLRsz8bNte4t36fM2C9lo/Y3GsDyqWlQtxpXVmKz9m7zRg20yvjKZrcu+T5dj
bB1b8SetstcCAiNS8kLxA14CF7HdBXvPpqysGuTXDmetuf5FTPVFfL9FFfe4fW2n
T7MqzDz7p6xQslj72j+AGMj3Rz7F1P7uL2bGqouq6hxr/aM0WPiUu3mYUwYjxwx0
leAC7FeLb+6rYNRzDQbqS1pukHr3asfUqkSbVvdL1Hy81pb+ndgv9bn+5xxXCL7e
2QkQ98/Cy1/WVo9V/zw7vjPNbNryaiDeTj+M/qi1qQG3dEScmRsuli8molL86YrI
UPEQcs5QL+UKUybsK1gu0mzZg/QK5YFgk8LrtdRSkpxA6vw8tDdUGJem8AGt3ssL
WQ1gUj1Xyq5ROQdtiw+qweHS2qOfSGitOS9WbpV2GZ9p8J4XMhVOUQinxuK2iJIY
wUR+pGSEEI4mOc1xiu9CABdsXkefgmz7YYqqhlTsHKcWfEbspB/M8JDS2tCgjIxr
Cxf/WGkOmOjBL/sfiAdwVdpDc46EKJV9Q2Fv0pwjL1RWEc+duQNgupfGwIkWSTaW
TuuXMI6zvGWNPiYPaMXYfGyU2Q98euBc3y8owcGXFev8YYoxDXBP3yKtmS56WyKb
Eu1F/G2dC10zd4HKw30+Hprt4ncE5SCbefbJYCZbRCaOoYxLsjLX8GDvoERJg1Av
XQfFDkLzmQWrJa/QVn8tPy3uFC0d+7bV933f/wSC3vSzSRaAierXGiR8dAU/bGl8
v9T2OJnS8bB6bzgIVvSFwg7ZLFGE72+8uX8CvUHNbik2URgdIzIod7p4poGd2IVg
lzITDNCeN+hJMZtSvkgFwkRzbGDzEW/NHAKSRxNrScugIwW+9YpqU04S6iykwJGw
7b5TeBEEkpGK6cylAHSBFNPGRssVi39PkPRXuIUh/73c7uW4z7G2YGrz335Yr/AL
n9VOjeTJnytq8lPUxJTX6UgbJriYtipTGcpbM26aROOOe6nHd1jcGeSxQ3rE8NbD
bohivHhv8GsewqDELDvSjpQ/Cy1AOrWw6GlQC5AQdbMIXuFOzgmgbyCybMs8nT7e
1Rqo5lCPNZ6ICP5qmCMK5fnPq//qCmLH5l6P783QOcpxI3uCQDREv0Jb8oMjL+I6
IGZ/tkxBAcW8XRIhi7qT99EphYXpVUUtwCkIxA2H9vIokdMZEPuMeZPKCleeCRSQ
IEisUq0gqXtQO0ckIsSaW0ZJVXMWD1cQ32Ro/RIpqAAly5QYbboTmCuvmRmFz+0H
YbUzfcaM1k7MEUl6KVgdxa+lAfQHalLc4UYlpSoUkvOj7/poSaTVT5NZbzhtPsaf
ZkztiaytNYkeOQ8VgsmSbR5XH1i6UEi0boEfx6wepdDPICpyKXmgDc+l9icIyc9G
Skimd+QiH/ZdZ3CPHkD/EyVc+h7XtKS5qWvVvOxy+m/1KB5H9LCr9WceRsC73SJX
89js6fpcMarUljxz5qRYqruLwCPVD2gJK53X1UysJgvUh/OTtoEe3fHRxXffkhR/
k7Cg0GopauYNplTCI9fzfZQXFU32GoVX+LCVv6gpKk14XY+HNObRe1UMwkOSdd9z
K52XxWNok9uz1gLVyl7L9KnhQ+/Bg4CWYRIo5ZU0CDmwVUBl/FVq3Lm9IvX7iG62
GilPL606WGWrCqn5JoJnuUQrZXy081ZrEcbdNyVu0sVDgey8Q9RWC1ZyoeMjCz88
ra8lCObdYDj4sTTaAEq8jOzHRBDvpUf3MZXRSVvwgGvfGvefHUJX6KXAgYeaiA+G
/vF2rCaMrCtT05wHe1fvhM2WXZ1N9aHXNZ8huVTaCwmyQaY5hhM5boRfR8WkJw+S
Yy60psVUclOnXtLPDubL5QsKUDZgZC2CY8YCnUHCYdO0li15itSik4LZrRrjiZbv
hf8F5A+GLgiY37ZWeATzIq5FgIjJKt0J31jns1W7gENw8z+N4g6i5Jm/nBBG6DN3
yv2Vi0ascFbdCNef698pyZFZt3jqbHRUbNA1tYGnTUQLxs7446zbu6fQ0AvNl99F
wArRP9oVCUJCgA9vihZspGAxU1QdsWHh8TzT7AEQjrL8YLOvYTaFvLMW0e1zFMiC
+5h6dY0i07gL2XksullwTla0RykqQSpqiVv7FEVi8LFccHQVVdU411JmIBwjd6/g
hA02fV+hWkwDcobLDyoYAWihyFArjLaF9BwT1+DXdbiWX/AzWF09k8PAqeAWhHwk
4T2bgSRwKmrdHJquwfW0zn/w/dyYJOZNpedfa+exWzgbOHZjhKhuupYTSpzwCHcu
ycoOA6Hoe0u0iVsibLI7L3joVwsJZzcSX6UjPtpxsXgmXMiniQ4i0Zp6cU1Z7idW
bdGH2zx1lzoF5bBhzsDuB+OF1aDCIfyZf4I5tYRbqWD9xB0Q0A4wK1lKvGeowDL2
PEQtFU3LzTaa5qpzlhLWAxV886jkj2D8ysbTcSWU2eWMbsc/lhgT4u8gf9ZLnuso
pVib9quXRCumFYL7uRMHbP+AKPcHSv4Q/28QGna+cV698nyogfcfhlEaNq1vahes
NOcgOCjRZWkkVm+ZavT3ezRHDMgKROHYGmQttrAS6Zahe/eI5sxDq4TAuJWhvoUj
lGPCgrn3ckDVL1uiC+hzbGfqPzN1Cn7trWpXesGF5qTPKmrVgAUrfhUJgjX2a5dE
KKNQ4gpwGZWuuJSnIiRO0en2uLKnP5dBvhA8I8y2KoeHcfWnj0ApxWKkbMtP+70T
sIHo6hkPNgekliPGhCHT+1pBJwJRkIGq0x/he8xoPYUvQQCxGN06XEpgBBk7+hxa
Sq+FdVCFbm5tQH0u0FxUJgykykPHmZjqVxyVwzsprXJn/zFiTo7xsgZD6Dl2UWVt
QpxIwga+YDzdzcizaDgvnQSHZz2JB+VhstBhL0TsuzkwGs7IKYepP0qNPYJ4RbXp
6LjnbPZsRbdDuIKkpnXwq+UCXtKP2pxxUMYGfraH0cfZMe6+D4nE4RivKsZwvMp/
T5fERSv+lHWsXNafc8fhUmdQKAyBrUEnTWNqgtc/ZQ2CHykx6GnULB5fuHII174f
70q3dMn7p7rfvK8a0EH/XK0NUlpQLZ6OKW+57z1u5a73UxMts12dGwt+fbi+QW1j
I0xORXTGfb89NB3cg2Uf02O2rLcyoaUnHWPbdMhLAuS5hxqi8Fs9PfvdiVnBHwWd
kM+ZhVYYfPP8AJC3eKJV0mvgEDEfaf13s5Tin/2cQ4ZQYz0IWizK4LjCiIerfk28
1r/6hZJR1YqjlSxVnVU3AUWdvlVMyyAceEoaY7yEMlS6tgXQkCHLcfkAZO/cw+Zb
EBTLfW49/iV3OrrtwDxqJPpK7wJjrQ3GDlddyaSIRDP057svokf9XVwiRJfFTa4x
Didkuh5IwUjPo7z9WaDC24In4Y7ioebzQOANjA2XQnkwJQKUTGyxjYwKns88sRL0
wMr+z5s7T6iYPv9251VJyLezGD5HXY/5YS/QdbPXnPMitY9kBQNUo5Y2J6minZDj
nIGL+AcfGsgLvgm3DBvW/XeLGW5HfMrmSGxoB1Us/4DRJBnG9O9NE1iTyCThLZCJ
TR92g5pIIXeVjw2zC1+Tpt6WEVDfg0qFkQDqOHMEzweDOK7zAqZtVPrjhz+/SXlL
U85xhvaGrK2P+Vtcp9DlEU1Y94n8c5xKJZXkTcOquC6E+BLYDO0/0UYulnAvBlGA
MFC1JqqnOjxfcY3JyTblUcQr6zzJOIQlrrU109fcqW5KEgJVuYi3TbixkS4yp9MA
RZZssF36MHU/IPmYXAqV+cST4hEtyX9watXqhe8+EebYVEZ/TxZWfEPNZpTW7f6H
1gJVPjObjeNqq39Sop6wawYtykPz2vW3ZzikYpcIyMQzhBk3WQ2Yv4nNao/3QvMo
1dVFIrj14I3VBQ/wRXriH4qcNBNNvyhvQsE7JBoAn9hecIne3RPI++HFHqnISu8h
Njud3pJRCUk03oTL1shGL5cmOyjqnitd58vIej/KVSQ4ZhTzVoSsmg38O+///4RK
IpEs+fE/TPqEMlz73qDPD+l7rbtTCxDb5jMIBNHQpNjM4Z0+ceFT219UMtOtrmyF
t6jSlXRVophwSxR6rLI1IvDhGHmKqJPez4FPmXFV/hKSlZxdPdepA4412qUvVF4p
hh6aYfCDPvfEZ/C2gXqgfgnm/jFMjEd6O6Ep1o7d9vf1a06gldZHfST4CLB/839H
c5wyVQvFSHt+S/k+TH8ge/NKlcYkfOZceP67GUplKHIpVE6TU0GMMOeHALxbmQvC
YrU2qLT08SWSnDWAc2il/+4+3a+Zc+tVZxgNAwHJH8gbvIofgHfWrHXejwjlr/2S
QujAzTbCvyxbYHNvp+FsCIea0GP4i95Ic6STKjWkUq94tq682ML74ZC2fu6jRqeU
7n7uu8qmVFvFWAZ6z18So6/bRrq2JqM0sKjy59wI6jXqkxGj43Azj0SgbrBf1bFv
5bhZHh1G0CktzgDdpPakjNO7uBGfePSnuu89BgNYdUvyK9/3GgrUinlUFGoNoqAs
u/eEEQnr3jPqrLpabMX8W+aWqX1lJRv9e00/sDmYPA+gB3Z3Z3k7o8Pt3diZ5U9r
BtEHPk7xJiouRXDj1HuCuz+S98ledu9eZly0SSFfJw4BKsq+8q2wAIUwObngmieL
uE85TARkDMK9UHb59cew+pF2csMl4d5rGqJjt8eAl07mrqBHlN4JKA6tsgBIAsqV
+1yhGMYd7gNUi1LLG6Jg3tqljVKRDIYGso0DhiBNg5kp93Zl3GBRIOrZ/Osn31VM
6A7wh4amReWD6htio+PmhzdZO0MxovyQKI33jOe6vIdGJVTqdPlV1YO9w+rHm468
F7sjSlRByw44gLjaJS2m9CUqi6J3JBSkGptea/U6BQYyHvAziz6yeh1sNOlFMWiq
joThT0Fmxw+ClzPWlCeKTyuJean9HCUp6J52w474zxBxE/NaE9kJH7wjMteXQqlE
Yyrd0Y9GjsVcqgz9igUBbLtY4WGqNZYSRREe5aghEnDQxGkZPfiN7huCBN8MXpZe
Ah50F9CJ0/zQzAJtcpfbuxxL2wOBfPnI5zN8zmF3bvVRoXjJNMLyeAhciXsas2W6
HmO0PLCiaFgotGvY6lbGRUgg1LP4TNmaGCjsIiHVvqm9ToGtcFRujI27IJJcu9AR
EgmutudCew03VHTQxTQP4aupry7/5cZymE9dpQYlzrt68pBF+EB9wSL20fmnlAB7
i8epm6+BfWDaYRqoIx+OWDQReYjacJ28H/U5va5vg66RjsOj19g8KMo9JlyJOH/8
ROVIvbQ0zg6K+qdzpA2tFhp0yKAtOFU05jIqppfubLifVXxVJ4GK3ctEZS6b2Qh4
4vJ/VBPhRaPjpEjNS0xuTrF0LpxxcBxK9i51I4/nTQQGOCm01P1mkUaBvn7ZPX+R
LiEGCZIUFt3DdkxDzWwGG/lAJgdviA5+vBiCJ3qe8QzxndaXpKeuHa1SLCdVQe3A
sH/oe+ike4hHvO6IYNcjzf75zQwqbgxPkJ0JHWVSzyyCIF0ghIuZqTZmWjmukXnC
k/Xf3/YmszAiuOMEKTP7SSiGAkNngHuxcViLhraUFAR1AU1o8+jqkZeL5DYo9VB3
yotEINwGGRh1/Aoch7alodBfdObuLJJyM21pO/XYpF2pKX9u1QvpohcRN5SG2XZ4
ndl3xHpf91NZxmSzCeTqhbAHTH7pT2ZhLAyzjPhsOuOzjmjhnuciIQMlcJcnaeQQ
/I132vl4c1//dj6Pw12tlPxAHa+OM4rdeXXN+SKDXxt+5mS9bmklMs4/wpUAfCq3
0UUya6Vqq96QsjUsCrCJo7KAy36X/D/o1/RWmFTuxGTL+YKdzKxt8gbKe0NINjrB
UtbXYVcZKAxImcvkkHVE4RvW9JknUnTdBpR2NiSepjV3tXwxV/TFAitBEbRa6YYk
a5gOFTqSI6SWNbReWcTvQ+DHpy/0XueAWQi4fOp3D6T6Us+gBvyWWeQGeeGUWBDV
gGxIHJ63yCObqYQgPJtZHs4aXvIhsncMhLQVK134buwJ9rqFaMr4sZabAeV0ZGBT
0f+ujy1w0NOQGvpOVhMVoiXfBOAMogYrQWx3IzJ+C4Nu+7zOfG7ruo5uZbpu7uT2
Kk1gpAevgyWoc/a1RTqjWKib2DSbsM9bCt8sIB6qThxcdXTswj79sF/iadAARw7Z
GyWNn9/gT5hEqy24WjvXOOF+rJ9JErjjxppWzB+XoS0JhE7PDUBEfvcNeVvLbLvP
mVjTUWRyVoH4FtbG6yHd22/UfBXJLi7SvThCOQJzFRheu3GCpvwiz5dpvuP2U+51
SBsSK6VED3jG7oN8yfyCRtL/qqcDDvZTTCS+Pu9nX0PB0ocANbz6CBLV6Ksq8AxE
y46SW31uv1oFkrDgTNUqFOcFC1QMmcjdU+bpfVlueSmI62K6f5/Qs/6WEjE84/Yb
RjXDMXjH5oXUFvrCa4EwP+hyDPHSX+svgRrs1JRkHzBIMdriMmIWcFcgvPHi+eXX
t5wdDw7AMtNvkaEzTiPyYY73kIvpEF6lnu9xXYbTY3TyEeHezH/CNmeoRlvmgu7j
NHdolOawsyllj5x53b/C7OtXsjcLKrlyw7fuihF77LYBhtahgnZCeMzrQ7N7FwM1
isuUn2+jY1Z6Rgb/ElUYxy8ha6nItm5w/PLaHBrE8wslaEmMGIO3ijx0Z6fPmNPk
T6iDHgl7EXyqhL+Ry6AH26b2qS+60MTii4fqCALXKKuTmik4D5G38UXy3gbWw2W5
O3JksZS19TDPeM94XyLb9eF+iSpVtP5zOg/s7nXRvNTfVYmTFyb08tmZoqi5eJCp
JTk8X19PeoSBiTsxss7gKR8Gw2u2hdyGmZ2p7YBIk6rPg2mdxOv9jfutVV9kZJv7
Fym5kfgYQ/n5hUQtEK5z3J604YTE0adpZAeJC9j1OYLpoHK5PJ8YT82b/bYBLKrV
HcIOz32A5TZkhCnEqUJWSvg4hxi+SGYqAmtB4Lr01AEmD1gV/IS2UXReUo8L4niJ
oOZm8grg0gM1wBJ8pEsEqIEsez3CpBo2FoV1scuHQmiFyYdI9h5eUSe1AhJXcwEM
eZ3R+gqDHGZt3+UrdShz0MDzRlcZre90shOlSGjyLYqaQOMtTh39UxU4bSZjRdJG
hT6whg7y2ziDF8OdPlIGQePxtV+84a1ZrzXCgAlVbSPNTiQv62PqRfHabG9+SpKw
JMl3xeOX4NzCp46QyaqVCCVGhRuadQW4fARzSjf12MYIplYXlQgfPkZIDUaXS5JS
iubmDP0/kqwfygk7oJ1lDhb+HFGzweAnwXbXEwgzbhI758p9cAE/yGWvSBtxuFxx
QcB0y/VS09WAxzcnBEU963k80KXh/maYftLDptjb0rzdw0miqNdcVPqhWsjvDecA
HgHRPlTMlVFAh0LpIaA/lpotH1Q7SQe7aH8wa0Ix7aW9URSPHPvjbox+vwKdEjqG
k9aPVLpBDHue+GwQ4UWrmsRGu6LDUTCNPHU/XiB/AZ0dp0smzyolF0uncAygMZIC
CYat46xe0AihVBKdny6IIgs9R0ltBY2aNqN/BFneezeWdubU6qz2MOcYsx2mY9do
UFxw/frLPVSiyqawaxrPvPEdFIGYhJc/uKsmAsdXTNRWc0gEJdaei29hmcCYbyMh
M3Ppui/7zBt2D1froBTxSgIQINnPW+5OsU8KulmOGAd0OoXkvGLtOo4qZX20nRRb
r3PIaXBcnzEBKUtkfjRRhsUjMgmDBudanB9stMV4zq6e0KIBNLhvHVOUne8ypx4z
YIRQapc6coAJB99yBg5OBGHEvzF7TTNVHdNx7Kl/xDdgD4bKj834GX5NlkTdmkdC
aB0ClqzUgvIruBStrXCFkbaWmEirmwN3OIYri1ia+CWr9EedZI+Ls7JWpaS0cQE6
i0nMnR7cKm/5pKHippF2IqmRsZ4iirHnarVyXNiiEqr2wJk1Z5vf6Nga2/lmAtUE
J2McViZH9n8I8yZwNLSb3k7HYSn1YBH8b2/D5hrsn2S5enJACVcjq1mugfFh1jXH
HnEMWYo9MBMYIs8HpBokmVgmPj8GFlQfvPW45+D0BUOnMK+7wBKdOvQ7ftkb95hi
Zzf6U4ljUT3TqsDj9upbyjg74ZVND9ItO32l4K2u1HJNh6P/IxGoZiNC/SSGpkLW
Z87XeOnUQ/UiG60c8oJt9yZpW1CNAVTvMfeeAlxZVTvwuMN2xISZ1ei+cq65qtMd
3npJmtRLPNWA+/lRWCvq/aiTl0sRAv+3KJZDEutixs2u7YlUxlreRNWvbhXjtNMJ
btSBE17vNoPnJcSiHAtlGFPB6KVnI2grEbDUC4I94hVC7BUhXRqGSrCrMmFa2Ors
yubtELDWfNcSxNyXmbReace/4hR5CsI57+jmB4Jy6sNzfMFD33EwdzjzyfIsH1lL
3z1E41QycSV1wyVeaVr7MzQGEwM4aDU1RqrbqduzMWJecemoMbjithpMTPtaVIcV
WuSe3XVuHtS21G0vNaG8uVRqNYcue0oMrNt1/OhzXV71T+yocZmxuYfYRmnkzv2z
KOE9e2ASo8tfsnaIK9bCFsXqkpxUIG2Og5PEZ+MDDjVadDfl7ubd/UpJR9bDYDDH
Zx4o1+QULaz9OCN25w45tsrTW+GGevJ0qQpMZhk4uG7NT1XkNPqhnlYFt+TPcapo
1nf5Jp0/W9S3RIzx9B7D8LH25F7r12Fgo9Qo/EcWvboDkA/uMRTtUKjaTCUhirwZ
oAZB3MRLLaRdf8xQA1c5+neEpmPMtJUc0dtvs5PvZmDbYP1/8oOp9akJIArLrk5R
czrsGmrzNYUX1iWFXiJBZUa9nST5of7FNZX/1c8ZT9akDYaDsUliy7ahtigAre3V
oOXSJdhReJbE2mHrQuQSAiqk0T4PF/HBl4v4QpXnVVmbbtp36olIM32sxQYVRNly
M4MGxHlcVEX1r94cEiKzmwIFycvOKTGNfsjUA2PDshXweZxNe6qcPYnd06loWuVZ
b2ZErLkRgnDKTfmCS58opOhIT3dEtnie+61XnSI2kznRGVlqqWIGEuIGQxOtrcIx
cLs+pmt0GbDW5e0Wp2VWyXagJY/I87//Nc2qntop2KbYQKTpNn5xVu+aH6nxlMtx
krVoy44hDJ8x6FXnC2MI5fjTehy1EEv5ZXoXtRfw3Xk+gRCQAL/Q0mJm0c0+9lZa
mGtnpp7B2MEvUCwpLPp/If9Cg5wnFtwaEczi6LIfMCc69G7WLwfdFcyum60KKbJl
6ueKY6qDBXzdBfgThhqP95xXwBfUlPtfRGisLwY5d9h8yh4XDB4Ha10hLYWl581w
ymeI8PtM52eXma5e5ul6jO0Vq46+jwtVM+Li1sPZHX5E5dAPz0cReGHBlujr0vTU
gr5uPg3zdHQKpaxmXLZuyFE0PNuHZVfBYSPLBAlvo8KarVaKfExTYsR521fBj0pd
8zetQfka5cuKi4GqvvvSIScf8/F6pJXiWI1CtNG+6BVk3wgQ0CqHSTo/iZ/HFEpD
Hm90wLUsnJPgQbdJryqUHvLTTWmhZ5qfRuB4DXeF6C8RC0WrESDvJi3ah6Nk/nwj
BB0i4mmJOz9tWI+ds9FgD58WNemEG7TNRD0qxa4/b3Yj6Q5R1HU+NuqfBI9dUsQF
QKBvb4xpI32H/6bgYZkwOvG9OnpEcqBxk07yyIO0xblhu+qtsqeFBop4xH04KBgC
OBNe1of3qetUkicDG0yyhxNresgfbNDKruq+s2a6WG0zCrjAo52x7b9Vdg967TrD
LoWkA810BC4BGuQpMvcMZPsBEMWxWjn1AhyFt2vGufg2Bf4T2Yv9bQTZ6sWlzCVu
lFmyYZU7seY+87EFsHE2bnDNanlWd+mLmv3OTNSJVolL2OJp31yr4qqeyKt2ss33
Gtu8RLkhhy3PjVtUOOve6SSPQrx6mc21GCeFLM/AUTU1KIigaKg48D9I+3XHV0jB
1KbvS4J2rEBoVzZbH4/jhOhQYAuz9AAESD4YmG7bVQF/Krq2ZW9lw3OI1cb2aAB1
979tbddgxTHoSfwmxBWxv7Gj9NtxUt/Zo3zmyP/1LR1/WD02NuIR9MqgKVMbsCFU
YQw2R6v0/Mql3G++mwq56uOLJjwb2k//O2Nht3Br3ErGgAGKO62DQtYvwg2q1Iz3
e+2lH0B0KaOa4tK8lS3+7oEuDLYuqWvsM9+PDTXqNlSliQHnzw0LpbPpm5rcR9DD
LxjnRziZDsPt4ZWTSeZURi8UV9ua4NhBbEunT/BZUrnJey65xu5+d6s43p/GrDAZ
NwLyVEN6U93R/2LJ+dzhx8n/YGaPfIpA0dYxtCAEkY921ctwn3NQn/tzm8T+vgIu
FKpLxhxInt9xnWvgPjshNELxLD3TUwHHW1v1E/hKgwVwD5DIbhUw5jXT9UfQGQrx
JnTG6OSueRrcSR6Pqqpl8uRzG0tjJqArScT35aogfkqCgZ9B9fDEm3bEEylIlS1m
E9EvVBrCou0DsxNeWPapjPKozTHTG/uAnWyTQoag+pdtc26VSdklBdLwPlzRVncD
Mw3HBwZvkxS+dbyAMt31Q4N1vGiGUH009FNSL4vJQhwMESKlXrtqAMUlog6Ccm/J
hO2bfmFny7g1FhhFiIU7TQNub1yB0M/W4FNbp1xrEGm2aIpOrdFbdwery3JfhRrI
MMTcGSPGXpVxLHjxYDDfdrG54pZXd38jmbXD1fHetY5NjRojbm44rurJQkt8OjAo
mDGmMlHdGFPo3+Aoagum+u7c2TYA9l8ejMsv8hzcrwS1kYZ9iFxye/JTRaG4Fosw
JYUps3EVrpstP82SgY/gMC5GGQaDb3QqVlTOdEum4iQPcmNL9pj+t/ERP9sqYnK4
Y2f3a0e4nWBcbOmN64PxTdqNEdNBJicq138b3hoS3NaYDIG8+hs/Yp0r5zZsZ9lu
OB4/W1llKSFpP6ZJcubxaQPtuVizm0T+KIAPKULifnlJ/rrjmE4QHjqdv646MZOF
PIMyIN2cQ/3XPj6n1xLno9duTn4BBQ1Iro6BJr4c9DbOUAl44IGeB0s/5lAG4VVs
w2LW8Um09niZvP3baQWfNA1fXr+FQVWmHw2Zg3mkCcMmLtxkSKMK5TjSYWCSw6c3
0PC/q4ryZkUf0L3AnKQgRUx4jRN8+WrvTBe0vnYCIasJm84qANPLWm9pNPkfcVO3
QIf3sbfpbYsKTPHLxNalH6iZnHUp/an1bM6rH1fn1PXZXlhipoyFykcpzPZMR08t
Psddvz97Rw+MouOvKiqmGkG8wsdrcKKLAJhbpTOsUK1XTE7IaBcEzoKcr7ja+XMB
R80mCrzXbWPuyGNRmljKKcb2s+JJLdNjObuGvpWgklsoHcNgBAf+JnaNpr7aE7zd
WW15keQ/JKuK3Ybtio9dx7J2oEhBZQ6p0wrORxCQaheEsjbdCUCBH1kt6Z+juENw
VYjpIWsBEudAC878XtJW1X3ssYdYdHr8C1F5oWKKbHXVXQ/9PMkTqziKJhskaI1B
qkzXXFOEVZvLnQqwhN4NGR5unTnClcGdtjKiqqCPAeghh6LB+aHswqa21r1twEqF
LMVdxTO86rfrxo9mk5dO78hMUBouDv7I4J/klLhkaxBlHAlCLIduqmFA6lhYW+hE
8lDn7dyW+r6mF4OMOz6qx1RfOu7XIcvyp9mapdOvW/AlHoIiTt1osrezZltzUx7X
/xnaRZEV0pST1PlfgJHLumw2OS5AzMzmbLUMPCjwlkRlLz8HIhtQxF3f44FzEY3l
AyAdUOq1BAL2r2sPw0dep6zBGwlkHJL44/4pdFWKqUbaZmOa8uaYKT6xDz8BRPAV
C1Zg9/ysBYLmQnZO9q/DXos4gmS2oakjnDkNxjl3ybibzSy/0a9aFWspjvYiiu6k
IjQwa3hFBBNvAOAL+obfPHavj70bqD77dxVNb+C5f9YsXQjnG2zTexXtBaXnx8ud
ogbm+BynvNouXyCKVi+7ZnTaDI/bZU+M9FXosHWWwJMcN+rQhkdXp9z6Q/IrZDB0
c33TXlT+q91zHRD4tFnRkBSVk+Ag5hv9MuUqLjf4zut19s+jvtDR7zN3pTG1KJNm
dUOhvk0YBoFnK4ChNm39Qu8PESG6jBlyEwd8P/VQC4Yqk5S1Px2ilC1qGRIFhbzl
/KSh9ph8vtmF7CkHq6VEp7S7EZD7radcb5WMrYoaCOvx0c9L52jhNJsE9zZCcsKI
lefkQO9heFBtAN+/JRMbwNjt023/rq+2jNCEq8bAQEKfFQF8k9R7kBv4a2y8HPIE
Iv/mG0KA7OqY6XazT2HkAxYmBP+koWMRotmYvrhydObQjqpdrUVhKN/PCVnAlcVx
+dgXW2PGcPUABE8e7MQliMwEbtLjbUzfx8esh7GsJkj/SjmsqaWohhVjJsPzS9Oe
4hyJSL6prTTnSmG+ztyqMyma7oJeTGh7xaHBu2oVXQUyobX501KdH+4r8LST3j1q
2zpFhn0AMFWg+yDOfKghZr9c92uDLFSYq+WkgE8dulcck2XUNVUgtwdR5pA0PQAy
e+v+1oV8NTsVgwnr5SVQkL8PFt/pQYi9fOVGdbN9rZquMuDkTya2mwYh8WA2PY82
PN7RLk+/1xbZuttIYns9JfC3+rq+U5HFFAWfPKENfFgGixcP48IWrw4wjyy4CBaU
3+S97vi73or8PJARi52jCnZqFBM2r9MnL0Rt+P+O4FIcwJ+Nnn92exw65v3rb5an
6+v49Zg04EYfM+/VLCbySllceDKqmWiUzjqU5n9LCsj/1SzVWKm9q0C6pueCutCd
XmBYTYBT8oW4/9vCrt4+/GxcOW4w56aYu3sISU/gmFHpvPxj4CM3L6z+fnZQ4lVJ
mxgtuk6og4Y3RxPV5exZwtXf/mvioKl0U7mVdj1Av+fDYVO0+2YgFbrxFq0Trfg7
NZ0pbv8TvheBpeCJJpffbE2ItzcDE8y4l2ZaOIfIPSXEaSxrcmRL3dx2myYjhMGK
HgihKm7KAVYwrheDcuj2LkyuhJMmZNQ1PRJB0hNKKQLB5PCUTZcKasf3j7QmU/nx
xKkJT26zVboS4woaRPxR8uO4491CB3/yaKrgPOoP/OkmcU5Up0XEtyPlovYuim8B
H5hc7AXkp5EDlNBnSWk48nP/8f1PvC+Her9ZI4oF0G3KcFtrEHZz3prS3fjLKW8p
NBZseAf1bi0ZxgZQeBlgKBRrS2d6MxQuSRA9+qYV8LLPcbZnml3N+dR2GcmpvMcl
R1fbvN4FP9T8cndTgJv/J4U7oyX7eDxF+HO/iNDspabz7sSrChPgapNgG97DbqMU
AytZ09l17inpn79zNjzIL02s0T9h8+0Ut67oTlvspbid6w97ygu2hOCGlE+4M3NR
iDrxEpj1QVcbcsO4eH+iqRgbQTo/hY7oHzIoUZD92RWaiGG62NGvpa3OHRaeM1CA
vo7EeMbEHik3FrmbuRND822ut9J5pPhDhalxdcR5qMYDKAJfEynedmZAzavCvpgi
xekbqWTuZ/f1RcRP1gdni/56VdKc8SKMNjzg6/UQ1Eqh2UEH0ABAnlM+ngxI/Dgu
xnzIEW+wH5tZxeCFh4Grfwzh1tzCOiv6yXZQyrJdltfv3xiuoD+d8s6yINvhQKUN
lJmzDOhSI5IpfsVl+06NSIwoq9YlaZEN43dZlzIYlqm2zZ9/8NJuxdBTrHzIpQmv
2vzZSAV0aGbypxdRboGkRQvP1/NbU0v0asaePnoWR1M+WLb0Ldia4saTIaOBdNzK
3HRP8xxLbsCZii8ZVCLnEwaZZGQUL6Ba5PvM4rK0OTvz421OnKdGFcglTlAMkx7C
a7eNq/kd5uXPOBOnmRAPskmRjDezkbP6g5o688hbaDe2152EJeQw4CUiVslPElzv
SlxUBaIUhs5AyiJdaM7/UnuxoRHRBp2u4nsf0JtZgJkCh0RHDW9bzGOSxuEfvb5a
5TXHx5POUg2t2an/Lg1/f/qu4rvxCp45PJSnnZz98WNQt9cqHll7ZIW4lDiKe5ua
n/T4rmj+x+IRVxVQse0LQgruCDLyPVgt6lkQ3wUujwP/Kat8Lhe1ThEx9zH0PCL+
Ox6Ywl4C2xD4cXUYiF76Lb3S9MMkzI0JW7uIKSGCeQJGrDtMzadrjPFTsJ1biQuT
shU7Pz2ubGKxX4FRl3w2IzvWKOUD+3gw7YRn51zSBxLbc7+E7sxEA04Xh2T00uzc
1NCIIwfTjtcJcoHY4kNWNEbv6vlmNord/nUz/o3EoOgUchEidfJWwmEqVQV3xaCj
19z9FED0TsHOjZY83BfpdgFR/wtQ827TMMEsgDhkkVKiYrFjgsWggcI0PliBVFYT
nbxI1Iq8tD0Ypsc+buDuecdfKM6J6oGU/qukt7KRuqCosOATYGwzfQEKygi3i29W
Hu7G+zIGkY0L1gPxDv9FvCJ/9/lDyuDHXseoMNk9V+7kWEDKU+zTi1xiQW2rnddM
MzvdeeyPakL/EMzXv2fFqlJvctZJ5qg6dHYQjE6TCXVoC2IDOi/ATWPo6s80uh8S
yeEbqnSqRozjOeYymtrp+gcvHTu6iYkS9ymUHixSi0FOCaCE0fHx6UhIUnp8zwcY
ta8iIiYjjLrR8MhE+Uex0u+M1h/CNwXl03v3QbpsMogAw3NWi8tyR6if4sAo8dch
HtN4tNIHAX1dLBtWpofhTzBntSXZkRXYZw9bcZFYwwHma3pC4ZBIvLIyDs0gRaRy
w6eO+icsavBsYanfJRlxjBKz1KxEtQrCT9fZSSY58gfJEfp2Q2+AjdiVwxe1Ri8c
3JD6Jv6EzKMfn5Ei/HmKRfoze+H0Gwkh95c2rTvG8WHpbfPHAV2h3iiMKeCOv32v
XEu4StqlJ6y2zFbA4qRv2zzMlXyWRWRmLMbXwm9PzzMM3Ezr3SAX1dpo8IYlgBa0
bF99h04WUXpLpyGYubH8UIjhlOYiQbmxxVd9d2LMZEe7IRoDvRvRkRWrhWURrkQM
bEfWee7L7E+onQzEkRreAvOT0XNCftueH+wcue6cRrFy/SXXRIdoMQhyqsXoyOZS
8IN1a9zRn07Xi1KPN1DUmwUNMufPwx2pZzil8kfhqIGSHI7n+pg0NlhvMsK65nRf
RGWgnHq82ihEOhrgcD0pu8o5fJ1N1Xo6niC0Get1vTj4UY+V5bFQq/EbUFp1RfgR
5W7qaIbtNrJ+S0odrtGXodV+4Yi7JapQKWz2gbR2KbmqwfQjSB5BVARb+NC2PiG4
JAknrrHkOODyh86w14mXzkD0GmR9YMjtgnLXY5aV9Kvrg+rfPUUqadx+O/EdepOG
YfoKS4KJL1HRhtiruN0PTWHCeV0yP6qFoi3DkkWR1ClLm3DqnsJ2zATTAslaJE6c
4NKh1fJ26Uir5zFIZ+FlmCsT4LKygl7lYOO3DIoyIh4v5YFcmNyg+ZuIDHV0eUUQ
VnKAiUhsLEwtpppnlOr+dbdXGRz7sAgD6agwHPdbBS4XQPHxEZMCUG5c4qX6ZY4Y
tlTtOAwuxCV4iEtwJQ+STfyiyCRNO3V5PJBUDzWqo4/583NEurWsZSL8r2aiQokK
5u24utMX4KB1DrKNeiTKt4WaCLKwvM8b2yruHTHblONnulx+ATkvFH0lKs+HaHNV
AA1l4+7ePBgqalXWw5z8U3FRfnvWZiBCPufO1hU7YDBKsni+GhxBK1H/X6zZvpkA
aqHOCobEp58WgqObnkbHGegcFdKjybCVdPSYyZBRTedKyCmCRvFL45ejZ8ib+zok
lUmgQMZ6qBtF5Z5p7lGyCwgYiBo7CndS5qlFf6MQb/C60gglNFkSgao88yk1rAyZ
/MinJl9KwgF2QDSNEERWTdRJZKovgC5xsNizGuB/V59unP6l8JHnZCkC7ejoUEhJ
lcQaXu6pS8/u9jsKjy7QRZ340R+DaP7GLU+fvswYMSeZmoqtgtqiwnK6lLjcqTko
Mbpn7JMOrzh/qJNWM3DJcTuGXTpTCoBMoYNS3r5ONDqOyQfRRJzYwxUKqNG+jSUR
o+wE3amu7BtQPctvztKxU8wwMz4+5qyfjVuJDxHPcfTi9Z0LCfEsSlSPFVPLxKNo
QYNg70RlpWxP2MxjCvskgcCaEQjM9raENqzOfPNDsCAg6ZLLo4EG88r/Dj3qtOrp
fF1EnTWJPH9yvNnq6a3CjX51XGfES2biJPBvcFjfLMXJDKwK9236vy86GzYQb+MX
pWoJgNoGelvRkXbF54Ytx3l0weYyKhEkcNBwQszmX88Jd5lcvMNUqQNekc9v5BvU
4Kq0mIIDu/iT1x/wphvjr5YEOgqdIprOqUBY6sH1N5sEokT40er57AgbpEQMRShf
vomhwxIJZlRAWnJn2XkU845luZFuq6IpzaSRQBgrW13G34Ja4vF4Sj/OPljVbRn+
8c32Vr1RVc5/BjYjkpCPK8Rf0kHhh+mxnkKVJUWt/mXWsMYSfVkzqWU6NRMxttib
XvPyWVkN881swRf7PzK06Tqw+qapxUo8fLopeBJVHeS0a9BIzGSqFGvWAIkt5Yrc
JjNqhnbd6Cr5qJCFg1VftfWHl7BpUxijIFpEOX4CRYeynBxlV7JQ3RI46iz2x6pw
4QRq9xrji+UCfRZJVwpFSRPlsQD6crTi4tDn0TiaghQwGlNByJhUlpmFkoMamUO+
Lb9k4e36aDznU608yxT8pD92i9vlqcU+pS8mTNRSbzk23+2o2mpDRDhLsYFrwnmT
ufGTgJp84cyo+SsAjSOhdPF2pdIAH5nEo5oIduOMFsuNUjNiloZ40BqX912ilpi1
VRnKJ9i0SAJfa6MZqSDuqvuVncpW2E6VSr3fTruvGwgohhaBFcKSb06lZZTXFxGJ
Apyrz8os7S7vQrn+jLAkgx/qATmQYpa45hMtFkScSFmKOCRcmsQU9ZgrXk6fq1eE
x7Xjbco/nvGW8nyCj7+xPjNPWOv/ayNLaJBWjdbbv14ZNEluwbpzUFxGix08/npQ
oT4t7ZHeZGALzCRBh5WoAKy96GTYftizq7PS751q1CRQfeP+Fji1PDzME+Q4eVeK
Dc5M3zL18w0EOx5mc3UH/rstChAK7M8qPRIiLcu4dLN/TxTxGHs3UFnyacEIKJb7
GQz93uZoK6q+gU3a0CY9a+s2JNUt+6a+9N1nwYj56IlTO9Abpu8wxbcwd3uxoz+Q
3jLY7ZPF3LqANkVErOXflVw/G+a/xOs8ebGetMt51/T1k0GS3aXN1+hJR9M8ZafB
oQQwO9dFbGprnLd7vjSnIYyJ+4/6T4pOaTISrlciBb6OJEcAjRdn1UE1eBGbkzvy
I+Eq4gFd7K8D+5pvXsE/heB+sT6xvPOAyRAhqfCCM2JFxM0Wpypk0nGR1RdEmPOF
tzZ1PkE5wz9MTc2Wi8BZK8RWHYnUl/FPaC4UnyBVgbzPyum7zNLOfYsoJDKvt/Vj
9Nlk3sPS2aX4h/YbJEJiO9it9TfZ/Ylc1dfaNrqCUlGrJgs1+AnmkTqL36FKSQ4w
pexvWtjmlnaAsOx7xKJ9ED/UzqHNVl+o/uBAYr2QUOytmrHRg6kQruUjFg7pnon7
T+62GeGILpp2De39LXoVydwNyopOQCAxagmitRadr7rJBmU64+HMI5RIM1PMujEL
q+1ZVaAf7gUuifbOVSJGEM8uBAMtgR3b7zil/iHvXTHo1mf2s4ayau8CromU/HCe
/uPA2rmXdswruSgWZ1bj3AUEEoM723GsROsn8RMeEGYD2mpnC3zKixtZHq3Jn99q
xaajekRXsgvCoRJaWNRSfEZgAXAigblKflrZVaBqh6y2bHtGgU7QGDuGcj/k2iRH
f2sStefAX8bVN8yd0ZKeoyKeep8Xan2GJcKDM042Ciq8rhOc2rFdfqQMZEnNVH/c
AECZH2vSu/MvfvZYDOSM5Rjg0XOiyVxCLe9gPAgdiDcl8cE6ub0x+HVQjM4KkzIU
pQ4u6g7gWY/WcU2Eyu2R82tllbF+GaXQ32GF/0wzyqubC5noWPuQCICZ/LnMfKej
eFSb/YHOIOwxdIsdiqOSHU59kpygqnqfCfmr3fwLt0kTnVS2PCSSNdvwaYX3CBjz
X11mCIGAtIUZQ03eWH1OER9X9BKizfJGGabTIxDH7nhvySl7sOKOrA73E4z86ymm
WxfwFRPIF/8ahn4f4s2e+jH/8BOfHvejOxhlQJ8XKvVfxOIb6tQJnQd94Q8irVRI
u26MNXGN9NWBIwzdY6fW/ILZqLLCOPfOVBe44dWwH6yJyOBkF8Uu/PKZ4KvEZ9AS
ySOGCE0pwJpYPv1/KHp0YUqTbPguXQBUOLe7CVZM9kpmgXAvBQtOmpqo1zLon9qh
7f0Y+SVA+woIn2a2pWVeYtnSotmylWbvgLADB0p/xLMu0Gdyo0jvd5drTMR3LbWd
wSdCQikV4dLryhIGxm7oJC2VzX3zWLxLZka+D+qNJs927tgfeJupOYpALbjGx2W8
/hCkO+dlrd0FF2s0592/+Du7V4u/F3R8eejPMIb6/hlHOpqHwzryCLeYLMdbUZsv
uJ7gWuC8vHEgLXCQ5f4gyR5UYi0OrjnSqArPmD6Swv2PVDTMzDpstJIwYiifH2hu
W9cpB2AdyvLcZsXiL5o91YbU4EcrUigoNUJpD4Iq+qrnqPLWNfAb0oYRNaBjlYDg
5dddvCAuqpOtG/jff4EeSbCAl2O76yOe7ywKil3Po/GO2MMxPeELN1tdVVstydPL
XJWFWvFcb82K01fKxSD6q4k+EJqSRMAUV+simJljrozra7uQub1BngUVhMZ3AT6b
vzTQ7i8EzMKcREnNWRwqPe+ln7ePStbnwJBHU81aBVtHTgJAMfJA2v7vEiTdns3P
E+L786zNn4N/pEWveXmHP8U0YH2jTYii0W0V6ssJFVwQxU/ucVN26RQrTJXTE4K7
KcdQclDo5Ymxs2Y6qH1R0lCLRn+WOzBuDLpJh1I9oYzWHmyNsDMtoQCHSd7lnlbp
xpG5IEJZeQfJL5MdhM2g+r0NK+++R326+ZJtdzc6TMXGlMEbexDtAR48+9gPgizG
omoMP023W+eNmI8nOvikOpsOJDWlXM1i/3IcYRdQzx+0i6qxVqgS8zhuDuGeyIm3
NHct1PVr3BpHy2rFfaOE0IgexQ9j1u4JbJQqTNgWfKCn/6uJHfyrVRn+Wne1u40o
R/lzUVCK5wGdusM3pifghlRtxuMPjnza+i40uBDDP1veUia5PQ0s3/6v6fwAOyyn
8E1zlJ5cUUE6695z0DfE8pbOAaks3Awzifn3ggA0sg/be+UpRum/+3hTiMx2bu6w
D3PuzEbNTtkR28V+wPj0PW7EOcpv4zDHk1ypFJN7bzOGN8YPvwcPMlCkI7gwMKeU
uBStGXzaUoU6HdO4GjyN8l2a1Xgn5UeS9twj4QlVuVLCNdcPHiOU0iAljXr+d6Bt
YTFKj9nIRdTenRkoHlBccmuToEHt0njXhn0tdoEOm/M04fJ78AWAIWDweGDglS62
ccdKDPbmIT4os4WUbICLkIlrpDQrQXsP/FPhfVeL+9ZAgxowO+x0IbjZzB9Fgmgh
qo3hU0jR6MbgwNXzbrMfA11DUXXN5dbTbNnPLwbRfmz9OkKvCMPz5tEKc2ZXeDNw
ryR6/tWu9F6X55qPkXQJIxq+RZeT5bD3qQlH7Koonbwv0jzFR9V6dOF6PD/uvleq
YGMvpQoBWG2J4YZLTkWbbRqfbSSxRgPHAQvx9AIzbmkhuX4lO1DRRV/LKYTst9Cv
O0Ll+gu34R6lpx+rnaN13VQ+BLjbHnTR51ZagXwH6GMm8zrFah32vQ6yvm4xVNol
tGQhWMWbfwsY5mZPDanH1uEyrwaV7GLtKlKJ9R6sXaegLXRDlDneUrkACR3nKBuG
qWlYet22cjfAvWXS5cChhyjL5gf10gmUFE4pw5ChwMWV3boZ9kgvLxNmKTPv7rEu
EittGcD/0dVbWtgUxtsgd3+CDwfN/K+PA3qPKjQDfkhwEo6/c5IOHFyidLoP7k3B
80iEMpENRlXQXA9fNrnkWEkCuFOJcVeW2tdVjbcsmckMFpPQbltaPvFLUVSBimw0
+Oyyz0LwuzvF3gnfTi7tltuLmjuMtZxEGH2L1srMo68ltGnJOaLND36wVn/K7RaM
D63gn45y9EbHqv8b6Ixonpqhcqr/2K8+mX3vcVrlN5f176qhG9eInRIINTpjjNnx
CW9UCAXahdGIsssZ5pHVweqJQlZHzl7B6ZLxzxjTYdemoI3vFOE2oF6J5jxfYEQc
SzlH7RGM+pDulALtK9WW3eDO31DNxxy7AoCuhaNk1MYgafJK/FCe4qwkeJhIDNvH
lgzsT91Cod6HfDKNv9ie0I9zO14OhAoUHcvmjhnXoa9xcG24xvyy/OPK4yPnC5PS
2MVenAFUhGEnvHsuH2uGZuS5yIDDEXcOuyCwLU+bAVfk22vDBpsqFwvsJZTNLGeR
duasfkI+/0mxuCGMpqUZJaitqxHMzMYc1Wk4RTi809xw63g42yU2fvvRLnxkKqV1
TZpZhMYF5muetdjtuBGunWtBP8M3Q2haicfP7hnBhFUBRo5u9PtmejII6+c0WvFZ
fbFy5z4t6mHDN0rLiosEaYqzbCXvI5YNBx1oH2iVH8ixr0nL4d4HHDFqR8wpGFdV
7WMO4tL6enrcIjJ2FNVoPsmlh7rk+ObT6TitqOarKD5T5PIN2uqUV6iQDC7FFMmx
6SbyiQwekqLbl6qVl6ibRI++TvAzGsMYHz+/x1O+Ym3M1kcKvcNDDyAdVbnKzeJv
R+m14jiutUci6RWQgAJLas5uAPWKu1eMXjs3rL/5Yg2wm2afNXPZoFLw3pvKs4GZ
RDTNe28/cxJrzkKZHIH41uVaKZzMPkdfQ/zn7qaL3SMuLX/3P6sSPaR0JnpSgjrT
r9mRUiY12zC2rWpIPQKGZzGneof7Ay+59tHCldMetkmRJtgwb41ny/6AhorLegWD
2lrHv3MxTFmJIYzVJy1czSMPX5j4Xe136a8LNs77pNQ51C1rW4FqiLsFRpEpXr3i
u10527WzzrqVJIENE4BXlh1FI6GOmkcFNYw/Up52cH6gmBvG1+/v6mEJWqVb0HG1
TUf9vIVUN8COUvpb9mDn5dfmgFK59Xv9l7D61U1egK0At9nWAbzdw3d3+2utYI+R
NTRAmZS9ILOC2vFO684hMhAJlyqOVKQ0fHq+0RvM0vjHvAcaIwT6/lVy3BGG2JxL
M2xRouprT9z0U2exm8+I4DSO0Du5RpEk9snLhJ4r/4pWVW4JBmS7bX//ZeAm7JIr
VohWSvmGQ29RtL5TxdteoDcuDUGG0AKdwKHg4JsnRSyAknveNTfnngq0WUrW55Gr
bgeZhsJ0DuEuZGcmS5wP8WASoFh45J9IVabSH75wVxGTg4rOPAqmgXQCrSXSncrl
JZcVrQ+Yr8w7FkrX/FTq/7Ml6XpAbHy9uaWcDua/dSP6YVfYlDcUyIiMC6iivM+E
ReXfV6EV1+cBnP/rRIqGD81rfdHhyJvkJ9enq3sbBmF57+fr5aF+ulAiX7Xwdrcn
uZCBwArwJ6zbiLeusoTFbekP7WakZzG1PVkESmBELhShLCfQXglOxnD6F2GjEY8w
S+m2qCI7Htn1zd80suHOBgh9eQypdrJ2/7BmlpniP7FSG4fFMV05VKr8a1Alsmb1
0Kj6/ooOoJj43+jIsbIG+C2WRcFP6Tt7XyvvhPCaKzGCoA1mCTU1kA94arYK6z6b
Hw0uPtWg/9dVRsTkgIJXEMxg7oZzID+WyWszPMkWQ/cu7SZJt8yOJGsxFbpFvjoi
0y7f5MDtij4dxBxYM09ME09WHT7wcIQO3FPHb8UM84Ni9CHPCFpN5l2bnCDZpM5H
r/Jj+jSV4eDwhrIWc3kwtXtNplKVS+wAhLUFhPcPOQpolEZ0EQgJBvdqdIATtHRX
KdmgGAwRHwE5uwBxgxSD3QvVRfaxOQ+0lAQDHEmJGd7+c2GcYlB6TnXb4a10BPz9
Mp8a8oeEq1bpyCgCJMdHdji66b8ZdfmMnF7PfkV1RBl/WO1EJl2qQnxdVbO9ZpnU
h/l/alrgI4keisPJMbMt+h7JuiVMDeNUxUUAHL9lK3FchUVuNo8Gd/hzM/pjRB1x
P746dsek85qlZFyadbUdrDPO4QUn94SAoFXALh0Knsp8mfa53AUUtmRVAD6cKmVj
k9kXsqPCNcRCUvyHsQ2xplz0WaxYVc6Ov47YRsLqXMYyzlQdmKTbdtKUdm5UnzZq
bPNTW1gRS00bd/MqtYaoqygHumDofGe4pVvb+JN4UDwggMGw3vIhf3e8wWhJsMSu
SO9OHHRkk5uVpkPUbOYRdACkImXPj++RawbvwlvIq4Sj/jXblbC51C850XOdA2BP
i1J0YwvZP4uKGt33IZtuABiW4PPJeYahhd3P1IJvtpQ4EDn5/0+RzUeo4Mz+XztZ
3G4DI9fAuMm7qKTWy/hk4fdwTABk7t0IytsGDfHrbHRVOqnN9IQWZdxI1MKtvWyf
7pjQ6KDAlRG6FZPy5bLsV/Rv5E8VC1+AUufrfroP5cho8arTJIP5Flhgot1vCB2D
lqALhNW+wmk+ip7G7Gw9Qo843qIDyVwaEyjaczy+tFshDaLIekvePUiU5F3V5iZ0
Pd6Mqe8VOLwV3mgmMh1aI+ywDP4fymIZ9VKe6pbNb7JmNQWD3TBlme4oVkOvdodl
KTvIepgg45SZpM4Z8VMufY/eRZvr2VgYhiqQgTMfbRIOndoEbfMxhm1IBQdcudVd
hm/WohzTGX9+qciU2BgeFJMhCKcbT+g12zdb4XZDQDaiT5dEUrZPG4U4NueqPr7U
WgcC0/PvdSf8loc4S9qWHj2WiSsq7CJAKJzQVRUYANhDb7k1h75ZmKJF1dsTSbK9
7igtO9efDs7MI9OQpR4rLfDF/Q+OjsUqlgzaPAyonWhVd2xJ+x4KZ36vKC4n+oua
CmTA05TRCn5POxGTihoVT4uqo8KlmphFDVc2kQg53aoULutt8W5YYX047irFU8xw
TxnZWFl07isOMD6ROe+weD06lpyauaGPCcjMREcFZgxuYAj5XSoQAglL2EzehJ5O
8AdPVPIEJogknFBdiMZL3e1eAOZhpAaXhGl2jIovdsgKbsewHdD4cYHk6tt8Qizl
GdDvv4r4pJotCr7A6BBvBgE5cBFeN81yDgi3HNFHX7lV8s0YVyCSzbNj4/7aF+hO
jEBZq+oyckgjkmJrR5OW/7xx2It2GERqgw33KAaWUJGIH3jYwuaQ0O1WfatkmqKy
oTIBpmOanKN9c2pe/mGhGpbdQh4SBmgPUvi5x+vJn5kOoyjOPlqhIHksAhKa4Twq
MlqBQdEl9ZgIXZPOzXPklKKM2Lu93jYOxMwuzzbdZkbKJTN8NlbihfGudlD/QPe3
06kXl+bzHTv5fIsMs+AxStyM8WfFuzUV/5ZTguaiU/nA0sGG3Dlss7IgEsu/ZAV0
/a/2ViiSDSPZMPKS43otuo/nK+l9sf1/5ldbstbx7Lcy5Y567mRcKMjSuiYHZoRn
Y+YdUxh5nXMAddej82nQEs4NXh2uZzenmpI7Z2Isru89yGgZVDerXQLhukwNPHb5
3Y0ZJebLvEz1Qrwdcqq6GC6stf90bzFQC9nYp0KN+Cd9LjCFPupCRJgxr8qWCiwJ
uN51f6ay1S7X5BGlRfWkryeuE8a0AUMMNCEashCy5JsPD7q2b/La9sTGBPHawnp+
dtOS1kVrCNauVPEuRJ7h8wqkp1cFkEmpNsGMc7IZw4jreeJcjAv64EJQEOnWAUFm
CuPgegbpiUxdpAsDfP+Uo148yLZ3aExrhGL8qJTNzougU/1sHev5+rJOBkNb1PP5
CCcGPXdxGExsa0ap3cyAiJRonJUQo+Flw89dpSc2nQieU9dWqQtajNSSs9K9829L
GY8C7g7uKGr6z2ZQIx+NVLU1BlkI8L2xa8dcL791oNH/qcKv/wQjEuOJXE5Jtb17
4qN/gmIiSPAIXGkBYexgU4AJwCYZKz2ntTLEDSjd3yFccvpbklla/vpeSApVhV/c
3Li1H9CdBy7YxE4Vsi4HT7MubJhBZXpI+/eMoRXPH2DBZ71E6R675BppHG5bz2Ia
t4Ou/YJc1t9KagqBmWDAOKZWIVCaoXuwuYULE3/HCK+7m9JWLTB1J4T3KaFUIDuM
TjwGc1tDQ+nsfZdGos/UrJA7hNSIkxiNSEnXnRPTCniaZQ6vPHY+tb6RXxP3fsfT
VPSN2g7U0BkNKhQSBTNadCxEeuTpGUWb672aOdEicOqEPWTcrugef5saEklSyD6S
GPeYmpJNBNqwXhY02S7ts27ifXwTKehsuSh/gIW+212rUfNF1+3VlijGNYuOTEa6
/r4F6nppi/Ht848huNxAWorilSlJLFQPvM7Qa948g49c4XqiOUcgd965pYcOJMCe
P+Eo4zTUsJKAWg79JIYstMGCWmlYXY4RpbzRx7jvxhteQI1Enbir+ZGCjkXZBGku
VF2cNrTHSbATyCcs4tJZiCvpkC86d2FtkxEqeFSdZmWYYc9vwNPlhbEOcA5zLJXs
BdDnoPmfb6DZAMdIO8xy72ru/ZxQD+LB4Z2+d9RpXkiHATL7GVSWXNHmfWR6IR/h
0n9jHDQfL/Rog6CiXKNbH9ygwpVSLnndw53m9YaKi0Isk9O07eEPEp8+aTg6YGKQ
fudv02wNNlnJh9RJCzquBhEWalinesQ5yIabGM3jJT28R7NgUt2LJRPBexruJSsN
1yK76vX3KKwbEZF62EFSedfw+LDIZO3qjzkBUon86q7DMFoOIEpPS2zX5X2cl2fn
sWnwOfp4jgMSGwuJutZfbHgpUdqjK+WXTElsbmSwSwKwnLzs2w6Y4uUGz1C8N7Eq
CEurGqDQWH0+6uiWL5LNsVZl65zmCNVJZKkkdSvuZEyyvvjp6QdpLwSuUTFXgyoc
qGueMut/CJjsCnVyRsUeV0/rSKo+ab45a81pBjD8UZ1XX3ZG6R4Qvj+rbafTg2gt
PXs3k7UrkH4TNwu7xFbJN3Kd+LHIT7pUt7/xoxiS3Tfu68JHV6ZObxYOxLnhKI2a
jg2LajWVMtGNXDfHfnlwxgFXcUUgke/06wxDwdlOfbHud24a71UgjnKoukafgNXc
Vs8HAfnp4yCO2eH5s9XXYoc3AWR1TkLG6ZDVednQjPj8vyzWDABHdeJmRL2flgik
BRw+84RwQxI32VO7iN+qnBTaKONp1O+3HpA/2AG356CEvVT1kNvGQDWUl4URKE1r
/6S+iUGkz+HxWS15LfjoUllss6EvarqIFm1vQ8iyEyebnSxLNETDLaIGGdQNFBtX
XnSIcnHyOE+YzmQMgyfa2zTdAk4ZWAr47B4bCbkLceIS/a/96JwJDExzk/vtDxgP
sKgFhhYvO9gehirsyTROZxIGfmsrOc+VryWwMLRqgIqA+abVRJiX6MATC+RWie1n
6aaGvFlQb+QqsEqirIs76dQLoMAJ7wPA7B2wfSIgu6QyOl6cLaPloGmDALxt0fLa
mR54LRM3RhhBdd4YgfCLyRMAV5eU9EW4Njnk4j4AtBShI3WsyL6+IEmjxYFNB5f6
NjRXI9saL4zQLaArgJJYIBVmWgYvwFSwGhNAeIHZiEjETtwr+DLYu95idywoodQF
EennlZ3ZIx1xPCvQ0/rfmI+pvMsG9/TZ9oaEdHjX+5eyvUu8e/TyIxUUNQTqyXi4
zayhZNcXbbjXAOCLY6alh2A1fIYwqf6vQc0RYVMyko/dIyAy5wnBFPg+/Bl0/1ia
E+mOMvUEmia+yIns5TzfiODj5k4LCpw870seSglQc/Kdu9R+puASfk19speKnPQE
UYw+ELgkGkn6szqYzUbr+u/kXuC2lVFhQ2EIhZjMfhagNo/AiyCDQSsSeC3AdYVJ
M+3BjBI8na/vvxTXp81vZg+lIFaSFY2BvFqaaZlqIJ5yMZ483dxMdQD9/6dXXAy6
2BtDNlljHxrsHMYdV89W8kErpHFekRWAnDkLCPKwgOP/DVpFZ9asiD7AMsQ98ldw
ynrtw/VePr/EKPJKUaQEBWBjK4WzMAGQvz8/kpZHStuTc1UBTRmhhmuDmLKCwgUo
3E9kqB40gwyZuOFhCtfV5/W11X+9pFYO+Q75CYWbucpvYUri4jbOcmPWd0QJGTdS
M37XP9U/joz6EFwK+EnzuyCSVJYVPj2sRCEOhS+iurvTyot6p8dYThgyD1KrM1AD
IECcR16dwPd6ZAH+cAvMSrInQmEgmEqEEcVAzTPkSxefXnhDx5E6l3akIU07/Tql
tEfVxZIow1j5pws6mmSOxoEvs8s9RobrvYP45go4ETJJ+iM2LRYbVaJM4yynQ9Xm
Yxj+X3clcsEniOdhcwxRVm5SPm/Gl9EK/9vetSTUJgShrFgP2Ge9jx3af3ahPAZ9
yKXumGLFeDuYb/zXFP2KVH4tW2Pm1VcArj5m3vI9E4NrzX1fJqlwMoHXpwEU/xMl
MuafgYebzTL84c+XAN/878PIl+Pd93azYB/otkolWiyaHE9f7FV5+AZCKVX7BkDD
QL2OyikYRqg1iD81GVA5imTeLfPe2/JkI5qkvhZYq0yl7ObafMQXfrHYGPMYTwkW
o2QDL1U5PCWJ1QNN0OV5O8SpN/DPk07OZxG0vAry8JADyrC04PNWuL406xuMq2QJ
juJfecwoDOfJFQBbnh4ef8qXZjrPgByj17XdTTzFqtALAQCFgSqOw0adUkRhae0P
PhD9hWAgiwwEOXnLzkk5z+9WIaXRbP8nTR7fy/8L/xbONPz8LevvmBEJFxHHFFu9
LyobutRawypdsn4/qXnsXV0GjgbCRF+9L9InjWvuL9G1pQvkf5/u+CApvEqPHd/g
4zrR8Xz4q/SaZvR4mmJpIFe+8xMFzte0XaI7+/GlBNd8l+nZEsYlwcOaaZnVPSvX
bGh1dwG/5xoElf1kCNC4r/GAuAc+6R/S+eGDkhCMMLwn2+viEpwe3JUc7VHU18Bd
aCEGuUVKHwbmA5V3DzIphRYnIN33F9/Zuu8tXao6GQq+kTDLXdXJxv/Kyo+mTOKY
+TpPbL+yRHruoKdukR5OEyV905umLY2TE7DCUVfGS5+lH1/wxWRNDkN//0/1lcgD
Awp3N9XiHgAKN2pFx23GU36atGlM3/d7ezXZKxJs5vS0K2ANuw/DiB0oF2GVlhWL
t04fz2cfe8UuLd7WOkUr6IuLCa9A9h9Yk051d0nN5M0ssMQYoqjg2X2Er86Ew9T2
GHlzpYKve8GM3olUF48ZeYy6vwn9LkodkB6AG30aLcln040miqiGaBrH6fSvc15r
UvSMQCUxXkQFCFS6R+FllqcludiE4LFqQUBIzbDgHo8vKza8iTZF0emYI90NFlOa
g2RRf0mxurXKyeLUXuQm8V9ewoAeiFS4znG+c8vi4s083z0c9qHtKPD4ZwcA5sJg
MPSBack8MyhWNHi2mgvOYZiZP8Fydsm8COAlHdD4MmrgSitv8lM5xvu7CwvJ3RRt
KMWesJM4v+HfTqWXxAWPVhdRZ0Duolua9Dphrd71DYtlmyHWiizfVseyl7D4NL79
moIzzutgxaQRiyKgTQ+dluyUZ5YAbDKX1zZLujIN1HKyAgB4Xbb+lGBBnjRKsM+X
sT5+KXOHaJkcviBheuhmSVQ1XxIzYJUznPSEtg8XVXDHjxRnBoNnR868FbV4yJjy
BB/Um1OamL4RPl6DldUYLDN7Uqcw3RJ7b3C5+sBdtCPeX+gxHNNiidE3JixyBpCk
ILVxWp3olYChGby8LU/UGjiAfMy2Y81FRFOd7ELV5ryOZtWQSs0U7QJYYe6ZRkFc
ol12C0t+z0g3NnphFlZycHkAI4EVFpQMQhZy8pY5wx3ov5d8LXsBp1idZVE+gDCq
rRZXNo/fL3wee+RcgNcA/P5fFd1iakYiCz9B4HMwA7JQX+cSaBTFHtRmTQlRHy5R
NjgnMKA9e9sDH3NSICULG+0hugwDLYDMzy7GiSW+DB0k1JsNwVL0GyPMWBtsibSw
+N4PS2l0E8zvj73GWj6ND1K0jDZavKVrhOETGoLLmZKHTew5yZpD97q8ll73YD32
qeKIaY+N6SFXXcrxosldRmZCYcp0aaA4e9+yIkU1NaCSmKmLS15vj9GdiGjf3uY4
ZGHphVjBeqYpIYn4HLhNL/+JJn11zyVmPm77Mkj+XhFXV8ANp78WlhOMvyW8bjzP
j2E/cW5Ve893dOA8FfF+GBhex1NxoqQEDGoLXeEqmDMYrq3AFj7niSfL0oTthyYW
bxIT7zIZTsyRUHkFy6BoibrD8ZDYl4qM1BySI96xXU71NKdPeA8cC+y+NLmdtFlm
uorBoCyTuqjtFYFgJFc4zC3rbZA8Bb0a4Wg6D2XyLeaE9FeoDNEX9SRDg8E6RZhW
meGMgup2GntsVXTDEqSwByBg4GmWLc/rCyjYkj0TK+p+UBDf1ftE2MMe48p8zp2/
xDJFgKV0oPh4gLnyXAZClzxaAO/4AuZ2M7YqnY0QWl3hK+4n469I+G5chBcRjUb5
8XoOSTg4m8ysngvUHSC4LFVWiTkQSvOZA59Q2z013WWW5Zb0J9HSnFprIU1wyYDp
jcbUq57xe/7RF99Qd0wcdxw9luMVkUi/3F2MnTsjwZT5IJqtJrcSTf8OydfTt9Vk
MYDmqbC40+UedqFQtpPt3nUd5TKJdHQCgd3Gci2Hz1cnK8JFAX8ojiu6aG3ktCG1
PFjuRWpflTXkBjzq4hXrwiXh2C+s3bv2+jg6efXYkaYqM3c3KuptqZ04Hapg6Wo+
zx2Unn6V+40TAM2scZX78ePdV7gxo2sZJjz7k6HtWZVVCB5NxUqYLOTeyzQn8OnZ
rg8p/kQQcc1zQ26xfBy+Qm072m1gVyhq+j5023pYUU9dtIEJZejna3FU5tcIHTZR
9XajDpsIoMy2nyLw3z8/p9J4kIkTn8LjUU/6rYwu4xT+Gbqhrwz6yfqQQotVOuK7
zFWT3StQe9W3WUkx2IpXvT9vV9oSl3YCdHgDI44bdeLPZULuOGXmazCfK4syCu+j
l/kNf5kiMxh2793XV4YIS1JHIernO8mDtSQpvVAM5e+VCZ2rYpzSbjiM6u8tu6RG
LOx9lYbep9D9OGy7jaZQSjccPaquHB2A6ci4zhYldvHFai/N260XGig1fPXPu2JP
RN0pnu1QXsPkW6LhE5pEV6LLdFC3lnuQS105ccZRpSUU17341X3SKT7E7o2UXVXj
yHj9VfSYmKQ71KjBe915sNBSyv/he6lc9cM4VFafkU7kGCoOShYcb61UIKY7Zinp
Bq+yZcrTkM9fwjlgeNyIiyP/sbdOuOol7DunHDUk9EPCryt0i7o54zbd0scyToW7
S2zoOJjlK52c56MnF1fQZtK3y2fTvdHiAxLCqKjavIOH/t5ETu2NWR53VtvUosbh
c7PZRxYqsPB8K7LgVZqrURuJz067nlPo53jlpTw1PEOqRLNf+Rx632o6rYtI//EF
AgPXXWAjBrqn23CL1N+BkZorO6ibU22tQtn74Ma07cGRhU+ziNCo0u+3IpB7oTU6
kwOYpZB53QM/djhCcNA6AgzzYWmKfyPJwfkCmzwMk0wle1GCJsPZJqmEO5N1vPkk
rWyNqOx3gU/WbTT2dNQrOu7xiXNHT+zJMo+mvjtxozrmQuFN6lPLu10EckVb1lGI
N/M2xhSuB9gzzPfQ9JD1v72XNrK5mLfZVWaBLDL0vWC4kHV/PjM+FezVrzAEShu1
U0NzK+I3DKzZpw0Y4fJCGHkBtWmKfmrwiPII6PtrHlOVyK17mvCoHzjkVTHpTxDZ
PW6S4djGQejzFSu4riuFo8YAvhtBzeyBNPX7VDmAN953sGSJHA/m/iOKFSEvSrr1
HN+8QSXq3RyQLyjp56SpwCQYTfJwCZjmVqfhFYwnI3+XFrBWxSmLDM1oDSF8a4ao
ZTwfebHP7SLEQPeyU8r1idsJJeijR+aWuXUmZ5uORcpMnRp4H7iDvwuo31JYX0B2
5jPRrOMHMT/1qoynZVyKFC+TeLqKxpgDhF+pysPg6FbdmpzewUx7HxQgK5p/kQIR
/HY8HwIMuaHCWnQf018EPF8CZNh9loH4tGPzNpYydNSzG/hBN6bTKdfuY54HHsHL
Qm990DItVWkhx0Q53pJptyXr/qrlX/QiKspY202p2xIfV3Ldtj2wfPULIqUkIv5q
dwpEzwCAOAvbFZ4C+mpJyLcz2rDbqXLO7EAylSqZqk0LetKtfY6mUMyb3Cc6dXtV
gsfVOG6nwpNdt57NrzmfQDdTlJzy7oFeahuTgNux1k8ydHNvse8iftW23YSg+cHE
Ks+bc9/AbX44ayIc3NYlxPSUwQZ/evAkMxsCeRj4vn97lfLn4I3AMxLGAs/mpz2q
kXqRDOwKqFsHnin0reBt2MVT3nHcndmRG+GGbleNCn4JzhcTHGo4MBvU7QjPzJqQ
3zuB/v6kwT0/KbckW1pxqDGaNdiFTDwB96ROcD1UoTC93cL0TgX1j74sf5lVfCa/
3KcjvSphh8tWVPd49SdrrGpHPaZzMsGuAS24tMhbGqp3AD8SerfDnHznoFOYZOxf
EcjxDdKBXY+psRqOZeIWarBy+S+PJXc19Se4U6nu2ehJzUfofvfd7FAeAewIP6Yx
3ifoBm2iaRdagzX6gOZL3c+LvouUTqvQj06FyF5YJH3mTW+r4PNlSHPHoJffo+LP
gI3QfOC7V7kmWcAWlZAfPZ/A6e+SY+8DR4mPQKcUZMnJ5N+pw12z1QsQREj1+tJs
FJhygj42O+rcOscKEPg6MnP8muCTDzC8wEWtwl6h1tDUB02eEYHxz13LhAExNbch
D1x/RiCJfvkrp9kqdupB9qSpb0e2YR454SgmhEhSXvWlZoDH+lizUfmuMIrzwZLg
2gM5yMbDOn2tmeAeMawc+1tAOeTsRtkfvzvKkZu0qZNt+l8V/7xukqluEnmfCGqc
k447Vr3L3c9pFGXFXXYUJqLQeH0UPSIYhzzAPuIUWkQAq2OmhCjastDkByonOZes
qoC3Zn6fbQaCIoijc0gh9DLXIF4kYiffcO9ni4IVV6vBqTETJ/cj2pMvqGng7Wu8
8Zk4hltYkIOPaef52QCRGYPs6GUSXrHzBvloLP9qS5llZvay3GLbmaRrn8GYYwjQ
6Mz7G7ThGiEC/HCTx0I9RFMChsdIjrV75jmFJo8oocS3K4CFKb4cRfVkjLnM2rD4
z/nl1HIGzf4V/XPlOIhpyG4cDD9fSseqD98HO/JAj/uD8K0tR22+sjFTwaLUOJJG
ZPupLLCwNG27pv6Com2gHeFc027MICzrhjCK9MpxndBXhMKwT0lr34Reu4uJMhb9
SXlKNGro4N2Mav21oW2emlf67JM78g4tSGhOlwwbxCsw/gC5sTUEQsGa0lPsp2fn
cwSGMVLbH77345bpHieZUMuPamFKpmg7z8d/nRXCp1El8XUapSqDc7iNFuQN6e4G
ahg1xiRN2GTzbefDvShSG9I7YemQOHPwAMMUYXtJrCptuDxcTmXO36WWx0Hib9te
W+MtVFjpZG/9/qFnc+5sR2w01mAsl0y63sN03ZJgAUgXumOUvAu6SamYFqG96zYy
1hIkygb8oIs1SiWNPcKZ/gZuVdPthwuso1HZV1+9e3By3r0SenIKqfNXK2Hr5/uq
c+voOmW+QuJVKyxUO0D60u0IeRNPYsEAE8pO1lz8NBeb8F/unx2TDvrEeT6DFFaR
evifdMIa5ZHq+/kzZe9mkQ5O1I09dteb3lRheikc6q1PT5eAUSBYYOgERI8z98i1
QvLHe/993aTGyCV1YbqfDK1jiMASQYZJwM1qezCTYYJsb7SJ76jhOOob+zWWj8/p
cnBlzY5kKwso+C9qCec6t9zVbH7RnY0eQs4trbJghERZu464JayFqLP6d2/PY5Z6
4vaJnLrv5fgF/U62D0VCpWMVmxpZZzKpFbPWsuLhsUGCYIS1ebwzQzfr8odyENhX
ZWyJGtSGJJ9M0a6DFjdF6zPpAyHdSfv3L29LekIAFpdzM6GSuhvDbABeUta0SVNn
GUepwa9o+KBmYWqBCyslCD2frLvMo0nUfr5sobweFbkMdiJX6XFhwkIi4lItSQme
GuxQWKW4eKL7LtkqDTbZy51KlHKMwbiYIfiBvqbrX6I64zlnfVrjoNE8F1nrZCL+
Lk75cLZGBFB8XRTzwZyg8rpDnn+QBVdfugyFArGxJMBpLP4No08HlMdl9y5bA0jR
jx5IjjEFv02cIA7FT/Dvf4VhemiX5AV/u8DBpykk0+s0L0uFMHcg0RpsP90swkhK
/8De/9wo6yEIuSCF73oLyMHuYQqwbrX8Uhd+0NngZ7o/LQDqxEFLVf+BQyOMdgWy
Z5Cgn0h2jagBJvKNpRqcEIxE/30+llXRbgkLZYgifhlpj9xP6SB1v3FLkrVKBrKX
FQseMem9Sjz8dIE8TOefD4mJ3Ph8lS0drHEPPb56B8JnDMSNXcXWvif3Axojg8Mc
eRiKy7HLpK15aInks8ukhJ00r9vhXwFHYFngL6xaTWJIW0yOH7xeKB8VjwELla/c
JmBDCXIvhithe6Q2KWv7ZooQFwWcObaZH+Jf+8/PvkRSO0JTrZzIYkeOhr4Flgcj
XGcpCmLcE8Tfih9SFwLpmDkIIOrK4P9Ugo271h/i0Bu4edm2GgtKiSPNkpZMFwpi
L+OrAfLQaqTT9EAOuAgUHiIdlOdZOf3ffjwg6crrFm95dxdVk+LWZ/ZuZ8qKQOpu
GA+V6Do7qo6SC3BTfiV2eBQPZawKwjCT7agBqU78RzWdm5GBjXQuEfOmN9EmdEtf
7oK8eMltKUGXxhBO/pPbj1glrvl/Ts81KmmBRnCHh8nZZRcogFuudBOoN+tBK7Rm
+F0IDudm1RlhZX3AJMBVr28C+cfKBYpHAMspKZREZbXhwBVj9unnY9eqHdTKepor
yzjbsRR3ZC+6oALrxKiOn/w/sUvM2PbOxPyesSFauq3QVGdYdKKOKUERMATBmDue
dMt5wZI/olxzRCa+5yBy8SEMO/e+MurIDkBdaxrv8KcOiC5z+aUSTBuz2wukccml
YNmGvD2rjJkaDABF3NWSe5vIkbSPCyj5yr4+sw0FPa9D/4xrzYtqU50PfCApEcdP
fSKabOrnjpxnNy6A1uVhpV9HyZ8a2bGNCQqt8Diz8wszwsnopcVAqDNNPuawkZwF
eKjHy4p/xOq7MHO3AzCjumfy6qe3nc7HAAy5N0wo2JGhZkZHGJ0YnjiHypa6M66x
IuDHT5lQaumWQeRdrRSmTCDLq57hwc9Z7HtVpOUEdvLB0sqX/uRBE9IL8a62JBe6
+4d2BHdRUeeQ+sKn6dGuSQxMDh0KMNvEVSljXQMGPbbQ8HuvdGvWs1mHf4gNEYhM
kIxBQURhV9xrZj6QJuw3PlKiq+jX0w/AUpQ1+OsSNLwrfrsoDKQ9untyBQRSNdhW
JlYd0v2U7nDTXbv4rY+jHBUgjKN0YdDqnNOO9LvR0jQNLrtNe3Qt72lj+ZGX1S2/
xN8HGg44nuzJ7cGja96mmly22Wmonj4vO2thub1tiuHI+XQr1iKGqVhoZS0Uu/TY
h3HqiFY0rJIXunSChM07N3u0rIEBB4bUcbbeVF6A/aNLbfkilj1C/p75PG4twwSM
cl5zvrLVBAqvx+S0B/vLmaBv35hfiE/UNUmBx+NK3jmvrfnEa3MJ8g+b95wuo9rW
vYyFVfN/78sGnpguR18tPPwnRkRQvHOSE7JVXBLlB4cXCOfbMrxudmMZrWO66YTs
Tda96tKjpyqropA1rtFU7+jWxREWG7hrEOElF/HqeMs1FzXJ115l86LItJKhcBRG
hXsVmbxPMWXWrqdE/tqnd70iByzVYHB2N/aDP0Yn0yuo2L3kJUf19AwNrtEEGw0d
B7e0Rl787RiyCJuEmtnSzimY1XW//CY4aGv5mb7xHjDhJO3BAqdh0ySjydlOYXvK
+lml1vpxN0Qn0TF2tJsHD1/I4/d0PbejHJ4gf44eJ2fqn1ybh7mNY08JsTqHnUYI
AJ06AsRuXvWCHTRSH4l3S3LfKx1eJ41Od4txs6tOu90W1A60BtNxyO8zxOvQVTVw
YiCkUF3HMK19Rcw4K7Qpa2nucuOA6fwFB7ZIzy6jMqtVt4gK+8rhfl5kjy14uWNh
1Of2yOjMPkiX8rB6n7iHfOTFewzphNDyGk+HupjnfHngTvdHdP94irpx4//K6lJq
eQvYU3SlTahlrZMmQtTZV1eAAtVK2A2c+XBzcY5xgkg2VgPK9QLZCcrksJGT5ks9
A9NSsjBnnsCa0h3wGGm8m3dYvRxEtLZHz/FYBSMvStzVublEhTGaSoK9f3gRv5xt
tYKsJhfqpX1N5EEZE8MXHS7x5Hmscm/HhBZtD82Ut0rM113n2OnpNWLQylo7EQfy
TVuhUWwD0tXs2Lprs3epvCsE6xNSHDJux19t1J578wuk45/0ChIRQ4GG2/xYB1sp
0n8GKjR0mf+bVp4f+yXaCQaVK2bIfeqSz8JMJ2Ia3pESLYelncxMxRAYr1MFq5B4
2wAS3qXQ+VPYQ9wDWyBNt06GEqrwsLtBs/hugRfQIR/Yz+7Bx+2bm+Sff1XIsNRU
C6BlnoRVEiTvqtaQZjf6dXIBnrXwtVGe5cqCG7wpcMQMZN9Dq5DHfiMkxYCvyEc7
YQfz+dQgMKezLR9CQl/IU9mgknuvo2wWqZhYHmyvvoI5zgSZx3LvOuRtKLiRaJ5N
U9/aunvR5zG4kwkYJ2ixJIzcuRLNxP6qL6PsNTNELxCA/qFnVdYajqyoehQctSoI
ECElkNMvUnnCq8LiNQR/tT4UVhvTdup8X5d2sVD5FAn9CbrO2TtOTDlrYol+Pk/4
aSReOPiD113qR8EfKMzgpbf+cAZ2kr+/hZIt6rPJAG3QOr9fbfxci7eSmyju1SnG
EtapdEGSzfc2fIuQKYYgRSncaX2BqKeV2OuVpyj2CYZJsTnsPniQqKK+GvCODgql
PVgDzHONo0PX+wYitS2+FWNmpgjNyhqN2LY2OMvBJt9KJk3VELvxL4b8Md08XYEz
jjUX+/kqMD7rEn8Z/vlALEZDtDp9Nsqv/lKKYO2LdPtnlz94O1gko7/3Hp832ruS
UG1J4l5swoWvRrwmUByXLQ3v1jNOHmEQw2NKaUznfaXrThLM5Xy5lGcNXlMun6/p
gid/Y2O3taNK6QVKCo/jhqiVq6H80wcZCPpm1NOJA6AOAC95X+jLbmAiWn2Ul95d
YAvSJEpdflfNz0FsOsNJ9Qafj9SsUi8gHF6LdQ3Skiux/ETmYqoZa4KuFozToi7s
Vq/FZ8fS7irP8SUqulr+Kum+qMcu/B7cEril6tgvvwG+Xy9SIjziguft6tkBpVAJ
bivNbxGWcW43Ge3InAxVYP8pcUCT2y/iORZD8t2SHIS1zWLpzHiGc5S/sI/o4wul
+Z1FRe2s/mm6q+8lurBpsfS9zrC+iikkq6OF+Hl8YNBune5P6XWtkQSfcOkcdgAU
2bK0K9AyF4CH7TmcPBoAhaYrKuw/+m2hp5VdZWXMfqW7+S+oFd8bBC1aXo5uwEWR
OgEscpHJgbW9seSnLhSJDfhxB/ZZaPyIw7qtGumDpyIwPhTIRMMHIx5EskgDMaVf
Nmd22bJOGXHVVv9U2C2gAWhEjMs7iTuv00BhRFJIGmuv35geqAn8CRoClQCXcMaK
k5GrU5UKIaIR18zPimusuYSscG+zsCtjiVp1EWa196OcYnm0NI9HhYaohzwzokms
xTbsQMQTsp5TmToAIW3OD/nu/qJ9WEfkrrZKt0X/eSgn/6c2HxJDphSfDPr9JjMd
16pcB86eDj3gwXb8DRyB07aMpGktVP6Pf6FmLnL8IeFDay6RfoS+nJu1zShWoBik
RfPMSDD3ZGYXxv8EIMFYfIegKJYIa5BNesYYULIQxHgd8nuqfP0W9FIyAumeTJU5
wL7y4ZFCT5mMHnPEgymfNOQVoYNTo/98pHS5ZFM8UtTYpg9nhCyTPqIGU83uLWQO
uDihCbQwkGm126fgK3MI5xb2LM9Mo+lraC0vtGsiW8VK3JPlIO3eZachXphkFJgX
SESVLbqeS2T6m7OpYMVcDfYPISQ0zjJLysZHkvjIBgttIXLWHxiOayOYwPN6JuT3
LxFLCvIPcxP2zdJlYwa04BaVcjyRGyCAuRK1z/QgnAsJVJPlqcjgsLynVkP4Bu/7
HtPAhO8PcxIc3kfHO+9zIfhPFIidaMN1woyjXfHF50KSWK7Py2rP/+Tx7vsJdKHh
mkcHjpgS3/7aGGcyyPh5P0IOqAi4Qhs35jKGb4+xuYdta7F2QpRxR3UM87PgzD4w
jLAqsDMTwaU0YqOwLoyljRtuYlSNAbeF4dPrFDc1iJu5zsgTlMlfmPMqcMXcK0qh
wvp7GLSru6DRXmJY18+M7XGnHRSKWhCRrxFM+HpQZyCCjb3VryxOC19j//yQqyHt
TQLv5tGa9gibHklRofIwVCd50pabepNMY+5y8AZ9fcds0qlqXvCeaWeZuHVI17Vi
vDmySdoiUoUlPlfjWQdy7cG8pR/dDy35OoU32X5emaUa1Om+6af751do19io+mrX
P8C6y+pIpmj3xmC1yMK3LeNN3ugofxntU+azFb3b8ykNeX2siHSR/uI1gcOpvVJ+
OE7QDrbky8YHe5u9QjxbQ/e38QaukPdoG2aaKmd/caDLE9bMudtwvBddV9KJhS6c
PseiTyjLCTY1N4TIJAkKHDbCV8dAUYxqnENjROJtUPm/dcQ2JOGNwodwesa8n9t9
4wVRlWKv+f0TeNO4kR8qzysaa67lbd2AKoctua09crd3/p4LxxV0msYpPEuvN9Lx
cxt9IpORJ0+452ZNwh7v34/iqgVJ11oB428JI+czW0qG0aCUEs/uS6BcbVu7L5mz
6AYfmh2+ECTxP4jREu6gL5XfgNiVDWjjlGMYIPGzoRR77DiEGJ7fvls7MhQQSI4n
zfiKDKkoYNknRsaLyP9odqA5H29g271nx7Oxj0lC+TGIQupd0iIzDZ62PQQGpc3c
Zqw1qbdqQ13dD3wcDi2Fd0m7NxreHaQaON31t4eJFvsW3qdYfPw2oAdpnD5fGXAE
9k/YQUDQQA/U1EZJVuZiKewDSqJ+ub5uhZCNPKMCnZ1fZYXK+IYO212aeompCbv/
NbSSZudyBMFN4brOzVVYWWKT4unGjnio4M3lTNU2FE4KXlSrs1oXKyelyLzhpdhA
6DzVlpQp8tHN+oGk9kYXdaealRY/BOJ/gnTUzweN2ms706gL+OeNmlB/NPgT1ZcL
TB5T0xxDjWyFFVCvYRT2MIEBWGV08XQcejpsyEQ2aecc+fKVI7FTXWWEvd8ZwGka
EqoB6hJg0Dvq+MZQyoM18ygUjRDqNAP9J0sFh3wy8+gkjh+AczUxkSFWpTzaChno
+GWs0N5kNSjq8saCTScbKoUtulsSPWSntgHgZJWN/ez4mLfXF/rmpCOYl15Rwpjz
xdWEVfQz8NMUSdDECh4ee7TD9PltmIltZD6KZa0AdzQ9Ekc3Mtp2+v1GOIJ2acSj
0ijWYntz1xpXU4+HJbL+4Whb8Mgtd6oYQplAFZyLBCLnED/qtA1zbyDosbDBmO/S
Pcg0OJUWe6aVhcYoryYC+BUzbor4Doo+UtHtQW9nI5kGA0n4fXE/QW6bZGYRGM7K
KoCoagtT7NFBlhkZdx9j0xdaOnvskGaOrpz5tdXB6p/AyvK/ruskUWf/m6bmg3bz
nyDZBidElzlWY9v+atrU3wkqvy0TzqUKH+JoCjJP6gAIBfzE7RjpuHfkbp9tWG47
uTLIbnUz30GVwiE3zCMObmGYqUu5IBykId1WYGb9P3YHquwfsK6JlZWtIEryH99c
CjZEeWcrJR5EMsWfwj0aIVi0mF+y77WUXbiBnzslGywYPJUzqZ6upiZ/sJ+KOG3F
VcVCfyirK5BPrj2ILC0b0gyd54PjzC0+v+DHRbXy+cfH2XGYjw9VjrCRYrnkEi7+
1PPbJcdgoO3GLfKZ94yiDhe0aKAOi9wzEf1NBMX2+OWnExtcyzvP4Di+UGiUj2l5
UWD2NnQ+G8r6Zzb8dokFnKrqUfpBhBSJRnHsEBw628Uxx6hz7xPWTPgzrqlYtFP2
dpaBgnJR6eiMtVc6wIUZ1QLxsObvghuig66fPpdPOjopPPJamfoyYIi8xP4RU5b5
UzLnvq+dVpWOKzAUZ1SYLykRpEktccjUBNXHKc+Mh48wrbAh8a0oWxUC4ix2hOPs
heOPe6rYfAXZwXNKmyO0O8XZMpmXLsBukrUHe3O74CuC4u9hPBimpznlfn+dlD0u
Xz6YD4ZOZtXMhCp2beLIkPpptrn7krzRATMKcdDSJEvPG2v8c+EXRp9/HUvTsiL8
X+1zB3kAV4yHqoamPbW9Ctn2YWhwpqhAySO4IPGJoSTgir5TkHkkzxZfhKqdptbX
DLskuBt+53ktqOLBDi1/FClNrIuZ/sd0UqkS//OXaJ3WQBoEe8/4Xotckd0xVdwC
87nH4B7kOLj5oIovRLxmOfZJz1yTfuyFKh/GN/sLM/e+WCw2fll4j3Fljyd9XLGR
+B9JmPdQ3HSZJnvWsWJGmWtygf60aKBkLjNAzeZmtcsmOnwSCwj1NO7ZD3gsalQb
Prh6Yb5FXD8VlSp1R5SM9D2nVT2Qykr+XjOuy9vba8Gq85Yqs0V86IDpZchRQkpl
7/igLbzyF3/k1LhIQc3Bb1HH16RKdXIXF/lKud2FnO7uK8JblR6iCo1bZQpKIU7J
BQ99U+pz0kVPE0MO27Nsncpas5u71JFEXlytrwZoRbB9lWJLFmSDkJMzUob6+cc1
SiOsqEpUn/vVOOp0uLC9wmBX1SUglCXkRFokwxXnZx00TfbP1sPCKZamlMDyzCzd
3kufA7i17Ns7VCLueQPevCHJkGpsHGku3/QGM7JboEyqDTTI3WylPivcfImnCHKs
9oW8nYjP5cNigrhXMasqeLsIl3zbMlEO6V1m+U6BbmbTSrH1/KMbQKdTYFNPa/DV
qY1TlcMEeox3jj0+o1YKGS9S2htbNTnPtcCe7EEtI53mspnA6q9SHVdNK1ha60Gk
pcDIOABXEszsCPfx9KUMMyvV+IiYLoZpH62LBBWCUQa5+uFurS/4OP+t2gGnAkik
71OczW2sIiWAF1bL9WCEh+lIXs3L5vpgCcqLpRdSIgXTin3+9XvnVQPfmLzp2V8t
LileasXoROORFEBsO/TnNwJhP7drGCTcNcL0BsUFEt1gpvK3KjDp6ccGBXYyaAJ3
jOgt4p9UvinZIYRoYOz6IZibr0To12wzYcOkV5+h4XaJSzqkMcjEr0Z1iMlRQ2Hy
g6RYgmR7huh2kmyCiWXPOkFq1yXBKQ3p5344rbkIsUNQsm4NTTFTw/ESOllJEY4R
a4XEMFc/IPW3vy1eOdMkBm538lbichxiWK7sR0D6lzzNB3U2gQZU+qxo+WVAFzB/
E4urrK4yAiDLk4tFpHUjq3Y/u94EMYyOzocgzFpWVHrL4+nT/BGRAnnoqoQUk/Fs
g8FzGCH5QtkgrTk6vR/HtAFwcqsq7hy/aRqBo1bMOzVDiBINuudFhbI3umXxOpDU
oHKA/lFDVAC+9s08oQQIkFFumvSul/G3RudwWKPlnAT0DBOtOMIU6/IaR6l/Ed9Q
8cVpxx7pqjFz42lc7PJdu1doD67YiZib/eN6KuWleZ7S/404+ZU4pam9wun8kNHX
VUqBqIXspkyD76jLReaBiP2eHt5F3N+dpbbMwRJQ8LyfqnXeFledEltA9/R7jV2O
tlXnYuXMs2HLtUeLp4cbCgwOj1Jeq55IeAop0jE7T84wOOC2PWHU+sM9tFCpfopJ
1wq3Pe/kGT88izUbZGPPjbdhbzvX2o2mKOhVHW7JkG0piBanAc8RBPgY9hFOHIP2
Qf2JUXseQ9C0tc2+FpUrWSwkz6tcgRfWPnurwXEMXWLx1GMWCxoaA2WZl31kHitb
yywgwA2LwuJNRKx7Cwz9jNJ59IvdiceHQrmjhAQ7tdQy9bOg45Tup1RUgMWA5weX
IuH1d6R25wPnH7/QRZzzWQVUVp3D1PDUvXvXOYVoFtXdrHOIVPdoGSIOcXMzzb09
X4zZ3jnbeGl6Ui8FNpunNxEL36e+zVth9te+WCziOr/DenzK8Y/C+0qEty01hLMO
n/Kna0OmHozaibfGCYGd75v620J8X7aUyPKPWf8SPESv9XBo281D725983nbTj8p
yzFAx5Qu3K8qu79C1C7UZ2p23g2+zjowSiickmNt2aIOP0cZzbiBherR02EAz0W3
XxBi4MMe0BKrywq6lq3puSDo2njtztsTeQoolTpwc9ujdbXriJymYZXl/hZUjoi9
B+AZSnJtxrlVZxQqo5ZsYXE7XIb5bTN9pPOfKx2+8zrm06XggpW5fCgNRGQg22uB
y5jXNYTFTEgPC8oyu9Rnqlw/jzPjlZzGIJAx/bFw2tjlUfNVVwBvC67Pcp3sbxSi
rg/QJsezeWxNBGo5ao8rRHpWOUjUEs7x5J7IFmYBrVTsJRgbDUMMBTZD+AHRmwLN
dRTx4R69m1y14GN3dZo56aZUYIKnjTqld0udIVU9nAu5IIMXZBVylDL2qsGwk5yG
7XgGoDDr+MfaZnnOyfm8p363z3J1QUD3A0Lda501bXRSetemkj9bFI7huLTZVBI5
JQ+Bf9OEwPiMpdTEVKkk65zDHYnndL9wyzD56FMcfg2NS6cQKg8usTvgGi5vYY/n
d0Ifrdgp6PGSpi1jlkdc2klIO1teI4Xi6+6+f3V7iKmNd+TTfXaNcQr7yPbKu0sP
ZDHfQdMavCKXD5dlJXZJnWg14fH39skiOodYps+gEbjYkklQthYkFo8avTRW3Nxw
8qFUzacePCqeDbpeP4udw9pWj7bWtCiJdKbfAO9zh9cMcemhfbIcxUJiLs7yvgQb
Kv+uVKDipu17gGIf+Tl3n/EYmUl0K3UXLulyYNpQlFnW6XKRJlV18lB+A+aKRYJi
GHbWbg2QsWEvaMbo86nvD/fvC/+bePZAm0gecSBZw2wN70kn6RHnrnb9tc/y3Qx7
RGHBk1RzVuTYdj0YqkF3Ng2WEs2150G4s4nnRAOTaJDgSPHyE0V9lxH1rhsfk8ai
iWeceoKUtLxIYhIapp1Mk5D8FwmaIZUh4H08ow1Ykecbj/NMQkmimqM6hjT74MSo
uG8HQ+MPDte1X9C+hvbDH4ETHXpBnm5a9IX9VxcVW1bZQ4ngbEgkmdmfXXHf8SMn
pNSUFbD+doIJiUxj9Bd9ePMibQSgzey+03zfyqy+xElvDbRm4VPnFCxYXMmK9mwc
NP46+WQRFnc1BrQooRA+Yjs7Uh5PxiFa431ELdAq+I1ea0T8xKsyvabUwHyvAp7J
RBZVFb3Q02dCs4A5ZDTjPLPnFcPD3u41Zl2783T7Gojtgzd07700EtBBVVrFFFby
4s72qVO+W1VaAfbHF8OdQ1SzcbiqEdA26AuWhtPYU/6YAONfdUy9Dy2GGBzltYrR
OShgYp8/mMohpdQR5WnacnRyW/bBu/8AczUBNFi4p3c7CyRP3s61S57ceAl6++Hp
vPM2YOyXIy6umhBsmPB4Em/oq7A4UgFBCkl4KR/9KedJBk4G7SPxOxLH/xqBCCLn
8A710ImRQxfmQX1/rACERQ/g0zKp1vgCmtEvr8mmq0UrnLZ282n++PfRMCkEEX+K
KlUrSsbut1XCgrOhaPfliA5jR5amSQqZeAIkVOZsKT7FylHpuLip30Xm0qJ71Ncp
q51LzIfdMGh7QzdYrKTF2utyxtxXkFgXfeGfzfDls/HC6XQWEtCFW4bgkKfbb1uD
WNBcUZqrbiaUVQyu/jGjDsSA7tYemAnxQRbPcfrhT9brBqiN3KPHUL6ozK6CvKY9
UVP7+WBNIbk5ItEyqcEdbGygTKrYf6iQr7dhT/n0F73Xwr7LwVtpFKle02CxsmQS
8gKh9nWLiU13v0DONhzCfRGfZNpzn7Kb7UeF7fTJ31zcoZ9jskorYWUK82C2ugT6
EKByEwQUSt8UR+/1ldzphYmlpIE5B4I2hgBdbQDU6JR5Ua46EwklNLFxV7Dh0oWK
BKjKAHlG1svE770vHJrYI8L2FAxjAAZjz1dYggJL0j/3X3htNR5N/cBzEo6iZFnh
JOPERxt6bURpwWZAFujtbyxgImYAvjS1Rfibid88lmTZ8ZLpr5vyVWjyGt8UAoY5
35+NDa+tCVPNjO/+u/9NlbaS58ikub3HGsVkUq0ZIBqjrUnzn5ekWwNn5+0wgE7P
+8veVMJ7plD0CAfXljCSta4od7+fdc0GGjJPquJVAy+JMW892uhWu/j66WSpcEuy
/5W6UmeMP2rsBPABg82FtiBz4G1SZJKOLTVebM6LjgIIR0cxWAMBjPBmKuuqvGXt
oV6XU/1vaJb0sEik5pLqMK4/GNZAAbdn7sFVHZIyaznrh2BGkCagIVN8p+UdfwWM
VKiPTWfQNVrXUoKHL0q50AgyR6DDHpR6rdJLe7s+QXRg2j8tMQU1rQZ0UH9zEh3W
elw+jCG9iet5sz7wXVuhhOCPWGbAmYfIR1hVzc5UxyT+2hknAKyvfqb07QtV5BzW
8TAohLPjz74+AqTFOsdXpqR3Ktttz5xbsAWiHZGUJ6nhIN2+WizH6XU9hRx2lQE7
ANmlYgSQ7YkaMgJvYOqmA0PbevIidxMF3AlkgliP5JsqalM8OReej7mVCk8nghJg
p2cxshEuzloSUjxvnSby7xzfeVW5Zs0pRT2mhu3kU8Cg/rCOC+ah6AMrHR4HkPFR
N84tADv1DE3EaZzyaLsVrZtyDsFTZnYdnDmLFvSnFl2UChzVLL9cL0ZBW6VOaIhr
WyluCMyQIlUOxoukKxeYTrJvBfYDeByJbuVdoyIurinirefBwWu9FYCbo5fQqVJe
q0JZOez5mQM3TNcg8ovt7nfgNONd8DjCSsfUXJCTkUWudzJ5qCmKo3v0S5RaXyU0
MvSWO8NEdSeEBSooTvp5/jr/iOVj/aptDH5yGL4h0fhHtz341vUfCF0JYiLNaBK3
qp2s5ymLStFJpTtm1hrpdp8gBN8dJXfXjhyncmv/9LmTUP0jEwgmw1fglUnbWFMR
p3zl1mt6014o1et9xq7EvaRGi2Q5l8gAXtayDz4bxtxEkySy8k5j/beipkckb+jQ
vpNq6Lan+EaENOQb44bMJO79TawRIMYPfRq8JjynBynp7neqtASxvmy8yHrDbFWF
X8uBpKDDVOyx/SWaIw80EFlC09eSlUmWJGyyXkccuIJ61/6aJsyJIgew9VTeKKrI
m/DWljCrQl+ljlQKt+et90OJ63c4UtSYYEq6AM2VjJtv7f15KjN7X2uHayROFtGA
tUHi7OcPyPHRyPlUyJHWqs6S09KPPLKeNDvak0uYSJsq4LOXLedNLgvJdRC9v142
ZXXtXVTiEcIUuYjlb3A0KAx5p3da922loKjk5A4vCn4I2H/xA7JEuQTPgHXSVp3y
etoKEcURoxFHX0igr93ue2HrNonyjfxOqNtpk5Fyq9a8rvjJlGbkL9wo2q4fmIBJ
DqrwawdkCOXfevaPa121V4B4PYxjdA218dM0vVpw78AIqbT7GMQXrP+MI8b+MiKk
bL51NNr0TeIxjrA3kdGOxCUsJVogSmsDNhOL89RpZjoJaArRVvN+PJVFcEgZzngt
be+FmycaggDNQgIJ/VFKAJbo25pfnNDMIfiQBqv9AvW8Hsfmo8oFoTHy8paYN51O
8SKAs8shb/cXiiUF/kbdUEpY3WH6TWL1ZjTcGmn9VicTzB5g9O/FsDfHhCbeALeQ
Kx6zfsGRu7+y6/U2vLNPzqL5clpK8WVmIYLdSjW6qw28sh2hJHT6ogX17aQh/Szb
xE3uevcG1TtNoEvf2/0eut9pxs7zNvXym4bs+DnY5w43exB0k9BWU8+zg+CrMmK3
UFXoey1CskRRCH1fLFP8UOZFUHEEqgbcxZTduPPWnlRxQFIixpjlkV/yuhWInJk3
Tr6A5OdB09VJb8tejxBixkV+QMXF58uHe6QPiodno9anbF0c148tnrabx/FOGZcP
nYC8EKeTltbfC0t/fB31e3reqgmp+g5jKSL0tcwH6+0JSJfNWsCbsXBaLZOlPGx0
eBjAHqKLCdGAnJOw8UoOGKuPB10nJFlNDlM9yVhpGPJ3eHKH3hEa+O+T6eGmYsXW
Ysw2cmo8jQpUMfMAFLYk6w8wKGRKVZQQhVuW8OqB0/d0i8mbQTL5aXi/rAc+QkHd
/rNchMXNHVtXOy0NhpKIRYqKh5jerDiE9wA5xbCoACx/0nNGr+Z6md7RcM7bN3JT
9KYW4SKp80//igB0+YBD89goO+vRvYi/FuUoZLty0uS/PhhrfBVhjhV1w2Z35Kr7
sUINUWkeSK5P5Trd1/V1f8NLDZQIz41w6Mu60MNlrOFn4h/LxoYFi/J/QH9HKEom
iy6yCgCaWx6UT5tx2QfccyDOSUq6xdU+y5L7cXs2z2ZI/G0v/cRE98uYJ7EESiY8
ibPjFu6r7HtN1h9cCtHQZG3ePY/Do1Pw+AyFaeok0nYP2i3PMF9TvkVjXC6lmJ9d
DQ//bwpjXw9q+ggypEJM9PpieyHyUBTEEl5k8H9Nf5719CmPcsz5+0jgiU3Sx2JL
DK6zblHqj2omMgYbQhmR+nrELJAP4FGFaMsVip/jdN3mtkM7oh0PEMqcYqGQKz6r
Rp0n9oCV85W5zHo5+Wv3wRvAAlWn6rdMzELCQ1k3L6LA9H4dC7kFVhruGlbVr0/z
xNbE3nKnChuuVCcp+q0DMPwPKqPyC5PkG6cp3Yg8kI/xKpY70ghS1YkGzILTpAIJ
J9WNNIdifwyfMzPL3EcBsICDogM1hBCO4a50j62KsyoQGhjRGAVjx+LEdwpFaVqB
UFBMgyobqzkg+VbKTDjUBKURsmAgLWT0ceQ7cdT7ka0msc7iyKJ/Sm6uNZ1GP/rX
Ome+EEJLA22QLqpOKPrV6r898ROpxx3hMnqs7KEUqIZudIqPaAU9qlSqC2faC/L1
Uya2gfRSKszlzzwFAXDL/Uf34CPpLQJijKWDtdpYtbivgBa9u5PI6eFAA20WFU5n
XoLrxL5gDVLiZwKRkh+0kyMX99cE4DKp7ddPLWSKeRPUeffsmpnSMh9yXpHsRNA0
uqLK/zURSbb5o19eQRCWR1rxicfUk8X1aftBfUgpNn//zmtIIaV2B8WPKsW2CZBU
MFgj4dfu3J5u7znNtC0QSCktpDOQFphfaYomqyskE8CqrRdjuvwhBL8FhLkA/BEt
aKPSsmptBsF+cw+IAPMYVr1Yga207D9zjlj895pXXDCSqU0/mTnCOKnkNGIMiwhm
Z9366H/uWNnywcta++5rTyUYrogome98ZZXRhlEEMFevckzuECm/6Y6bh7PCyTXW
ZfdEds7niZWHGXrwRzy6VsFLkSCq4Z9acdyTXjb9eKurADYwl2iJYbqbu+CAW7jp
VF7m/EHhg/5jhpf/lifcNe4C/VW+jG8ep92m2CbrSyyhoXgP2fXFY/HMaIU5MaCC
XUOYF3OWX0lONAGqPye7G7aTzZrz56mIshVsl5U4EjEnddzdM9QyqTbn7CQKMCae
GxpeEcb6WEDWxxyhga+gRj8Ju8ESTw8RkGFDekbvga4zOMYOed5EzelwDlId0GAV
9TyPiHYfGbxtUygDgn79w0vfsEg4yQyhuD90PqXkFLuJElquUBTP1e9mnjMz1N+k
v7i8YJOg/hhqLQX0NIqJ7IHiMjWCL8RdtqI8qt2HncbS/lESs+jeXmzpSCg6Vu7y
OFHTJN3bUHC+IsDLwWJCtGN9FUimbemPlziS1CuRSh2VI3XOQz+UQPvG43LaCePu
ChnqGbEU8b5yfDyN9Q0xYwI4cz4GSVxJn35MhL/0Atvmw+GfwXYkQ3yhq1RjDcoh
VS8P5FU5UY16KC/JJBXlHRlr4/McFNUKM5KRKUEwTxJ/wAXb7JJ5ByR7vBjNIF1V
BKy5YwOSf33nb+aSii0ZL4KuBZvqAACzTJeJ9+R53Kz9k7XFih5lhSqo1vXGECC6
Q26Shelzg84LAUAYZWZjG2R5g0n2rgKs8FpVmAPEdbpSbUqz55drS+V4nMHIUHsg
4F9DCuz/uey5toSvB2360VahFU097Ex9G1mz7tsPX4mUqGuT+s86gvuB9PURG+ys
2P2rzVqMaYhhVTsz0YXBVnmBDXAGOs9lCY5coRVq96h78c3zdkOrrJDd2lumZS/f
c9UX6gqRarrjlVeMZEmaE/j5h439xnhZwyTtTLYp43myXKAEC8zWox3anCM9eqMI
C/JIg2RmLXNDWTsqU8hjptXq0Vctgb+LsfgqCU0f6XU+2v2KkMckcCHi08AL8une
6TDjp+rOeK920trTs3UzDX9i21Dv7PMD0kMdA/edfsOVwlwuNAIElQKibh64n88l
0i2ilH7PFaLfF2OYJC9f4o2gv6aA0Cb7u4bRHZ/Yfx+REv7va2eU0T/VnbsOF3kU
OV8eWwDmCCmglHi60YnyPPAG7eKkrod7rv9TobZR8NMj3cQRhZRBPAybyyx+GaQO
gYRjDyRli97jAx9ZOkz5beTv+THSkJRI0bhvHnMTouaqq3RnOtjuf9shVcu243bo
eFkSn581ir7WOj7ekt2YDhgs2ePHl+HTS60BTVx+PHitZsbBvmMUUMfYEJZZ1U2j
y+iwbIjuVEj+4jrod/JU+4J79LUbhFeIDXORLs5MzmZ8M8+Z9DIiyC68WENt+BJl
cUx1v9BHwCY//llRx3+OfIGHhSEtTEZOZyltp+wD+tPIuyJ4mrOd6m6bhQNXU733
xkNU5g2KAdPYX2bzWtu9bKoXbB5lqvv7/+x20X3PYl9wh67xXO06CFbhy8oz83/4
vxK1V48kezEdzK1zYuQb531fDNfzeLARMX1/ZsTaDEV72C1dQjVBfcDZO8pkMJQX
4sborXTBXxokcmHO09gKefyckcgKeFddgWPL+TmbS8+kTz0u0lHdlJuqfIEN1Qcd
JQTt6fVzj1TXY7+LFoJTkUn5e/xKpUz6sF7bLoWnNKajBob2sOrMoCHeX6vU39FH
ECCIqQ41FYR599vIYSYWoZRYBUDDuyERN65mfHR9kyiVusbj+N1tyJDAJUTxI2bb
fGYLQBDsnFqOnQ0fgjaxmyFcss5gQaV0E7Dw8SAGaY+JNsG7Ba5zBEoqVwSKZ5pb
zwt/heg5JCUdcPFQGyIEBerN9vfcovet2jB+e/UfLDYlrAta27g8NsaxqcF+Xy4l
4jA6whg6DOWHMMR1tAvQBAlrlLLZuQrwz35zeJRGUyLAKuf0uAuzCMfRe7LdDUEu
KorUNCtUVH5RHWTksIfEK1IcQMRj/QgPRGbblWVDBYDrghk1ZAF0KZQ/2R5lh7AR
xjWhXjmKUEK/Tdduy2dWE7ZZEmpV/108a2vc/1Ly6KQY19vTcMa0YLeTKPiwOuA7
/ikqD0Q/Ud1r8tahKUSiayYra38fFzUNy7aJNig90juCb+ZR7IH0C6isdR8Cyq+9
pFrwduE40eFpp1p9DF7WO6Ks3eUznGFzdtZeNUyOk92xxiVcl9lP9R44zckQPnUE
eM4kX6dgFUWokCKSGrroVj/ypDobLYAysd8+dAMK4iRL/WUsKElYD1dCuWrLfunI
cMuIhJce4UytdO4iINlIYWDflusfbVAHYOccUpMpQ+y8Iw3Ydb9WrR/wxHQ3Gv4p
excpJ09amCgpv0yqmZl8PBk70Jd/oJYjbdbLBRauOxFQvGZVKiN9PfpRWlgnKMVb
nBzgY3jxe/4l2tLg3GgNHdaqJEu9yZLVD0XElLDYHi3uTH3gi3X9RMTa+jq2eZaA
s3KlvqIWXH2h3JovX3/fnrx5LygoBdpnwr/JdQH2zWJulfDCN6MzuhhuGbFPllr0
4XkYzr7Zs9yK4LAUMl0nC/CFzxCfchIhPmyQqraYCv7WameCqFBNRQCmbKzso0iN
NdBZqEU6LqCVjvNJohPGtOF9yhAEmuAvYqpkUH9sRD5Diq3OoIHdkvBdtH19v30z
2ymnqU6FhQ625j5yQ5BBjEvsq8W+cEJG8OkXYoP+NtWBcU7cGP+G500hkdW+0Qzq
2kqDcsR99whvW7WUCaKlrtwZO2bnwGoyoNXlE0M/O6Mp/iCQT+5irqrc/HY5QSKN
BpGD8Kca6TLwxolXOMzntDc0pbvq2eoQ06sD4TDXvKOx+FsWIF1eivihv3CndBnU
m9V7j2leDnjQFSh1RmxJo+08a5mSwytW98RVlh3Kay+pwSdBGWTZoSQJ3LKBI5xM
PckxP7rrdlCDPXnfxkUzOn++5EsmtppQlBKIfsEoDkp2x1GOHc6ksndsQGP/kTla
O0y13H+yuPflY7tj19FJuEK8bAVkLjy5uDnkJiaMyNqklbjmDORjrbJ1E5IMyvvV
5xFEusybuI2tni73r9PDAuHBirKaaI2TFvZ5gXSCb6a1QANjbLIGegj+1CAKq4RW
qvk/cYTJyPQvJDj8El8leU8KGPFiHiYcUrOpF6KmvOK7PnvrhcS9mz6ZkP/wuBQV
47oFv2JNE3K0jR3qdPd5TNb95wp9aUvGV4C5Wk+2vsbRstYA7408x1pqSxNe0+5E
lB29S2IdlPcAhcSb+XZw017uGZk0BUF00B1rkc1GdkgeluzbUGMwgJ9GLljPF3q2
DzX4Pma4uUUIBa5ncyP3HGc/uJMnKWty6A5R8kPilSSCEg511tZxTaGoiuLhGInx
MQnHuWEPS1BTGTvjvM5aRfgZwmu5BF8WugO4F6c0IJtc6naGJ/+n94ZIaeA5F9zv
n5uPED5YOPdXOlb22Y5TTHucv+jVzBasKm34KnDokis5r8cZW6VEo2xYvlt9VSfb
WxNSkvdWMoSMtefRB47E5UqzX7qJTYnfypOztcT1ljW1YFP1VrVr8QlNx9YmlIxu
/b4DZIjulkoFBtri58P1PhIuORlP+1UIhxHZqV9NMqZQ67Ai/fheDAhT7UdSsHEq
CWKndtcOTFy/eQGwUJ5Kwp5fLvVUW/UMN3OV/SnoD9qazOeXE8leayC1JB/4yom9
Fq9sFDxtL8JfdhzFTtB1MXZDo7H1Rs5PHagICnzWhFNndE2yKrHA3kK7Mu95i5Nm
2/VrWMzoeUyh9h9zIpcG9JmZlOgbub1W7Yw4q49iG1jagJYOtCknQXxu0uEcedtk
b9Ph4MSEen8WxxmcrYG59majgGD5iT1dKm1+T7X0M+YvuNqBYpnwAOPTzddTZpjN
fcy76em5tW1RW9NEqX9oJcyO+Jd4eyi0zW6I5wfqpDbSQgLF4Xxt5a16FzcV73BH
QY5QfJKdQC6zeegXIdRATYi5NMFTuVacsYG3gQDkxVsR8ez3lJ+cFkfNMiJjfw+u
Ble6GvRNVSZEvUzYfMKhg7fW3ICqZGnjSLYKYvAfosEvNQeHBQ68+lnyfzBONRTc
dCRHQbp25UsXwUI12+iw4vTsa3pFtoaDHX/NF+zXO52EFSBlIaPHAWxEcnjoMPkk
rgfWuM48oBripgiq9rbUJLBKY0AcZmeVv4gu3mSB2egMTHHlIoH2gIz/7Xh5zn7y
nAkpeB4dsV81GrX5LuG7TduGXJm36oemsvCnhLmxgVOEJHkUd6wVVKAkp5nNMDEh
lUOgjhdhuCtoMz4yPdrYv7N58YMYigNDuPy4cwJFhPAg+NZ1w70mfd1zVltDn/NT
TyHu2fLYAXOx8WnmBgMcRr9lgXbHHzyypmJR79fazmPkXlxxkE5uHDyS+ji+GJCd
wbAVTczdL7+7hgqebQwKsmOzPW+3Rpnm32rh2j8BY5JNS8uv2RJUNFDuKqlrHiZO
wS3H3T3+L+6b+AzNnbANnyoqVKYd0GTqltprA6gH8CZakaT81AfQijsF5yFEgB1Y
AbTB3/MdaXe0Mp7Cmm00j1bCCUc8OEZffhsefE5ScDR+FahzCn36MwfPtNxMO4dH
hXeGrc/Qv5j39G1ugt1Ef6mMgXEXVNj4iSyCIbvu3vQg5Kb+uI97QdJKZeDyQrEZ
YWMbrfNjcS8vuW6qzy8R9xJuEGcOmbb4JRo9v8XZF1Phkb1sLKne8QMKJK84vd2p
LH/QIFQ8q08pEpxYJrRmftg5nXqypKqxKiiVcmtFd6CMnU6Wr2vuKfIBpp4Zc0Vc
NBbjv6kSHpq2AIiM00OCHt4L3cqAWvSdp5vJVDYbXmaHV3bdkfPjZ/uHhkFfWrpd
83rAc76ahBqr5CqvoHM8fp0CFXpiBeGRgliDUiSect+Ap5tcjgLrmywCeIM3LxI2
RHSK8UcC81oQeNhqZ58hn9bA6/OHgSa8jGGURDULUfCBzJNO5GqN5fOVg/PHS0u2
DrSTfoU1xiCugz300fLi0HOMM2nx8EMySHsUOLPfPfs8QPc5l1CUSX5DA/Kc0wIL
1EWfkBFEj48a0iJgxTU9ihid3JZ1bbBrByfIyGBJwOeA2h98DI+e0DB73wC0DQWd
C3osOiWWPRfM0ID4De5vEgY+dl4eMMMy2d/1KFGB9yQCWlUNihuaCUZoGrAkSDmy
3lAyylruXR9toHskaucFrqS1kgipd66N5b/P+ykHePx7Q7Q0L/EWYhkq7QnkLHTa
vd8+rfZM2BUlFUM50/OZo7ieCz6HPTULs3u1KGA9x+nK2cDjB+KiTR3a+WucD5v8
eXVo+Ae7f7B6OTwhd88zaT5l4bLEVqTexzLA/Ucz+hd7Uq5E0OTBLaYmWwanENTx
YEgJXIG89jMm7h/qivaNPqVect2PFz+pbZ4GbJYT1B7pYnmq9NYHX5/xBAmDhN/p
yOn5TdgsJYUoO6IXsAc0tQ3n/XK/bm2Si4kj8yiT7d372OFMZVgXOoTaSUaEH4gd
cWTEopevNPwM/TGu22q0+jIOuwE5HjilYHXewlW3AeC6h4JyQBRcdzbXrQpIr+yc
XQiEtCIP3iiqneHtdGcX9jinqwByK/O4AAeH+G3LCT6JkWGuJCZ43fsVNOrSgJva
OzHgGIOm9htkXxRIo2XVduq4+pLBEYGDU3fQlD+4mO7nsunsOYpdco5KcZ782AlF
5i0Mr7XFfHoeTlzpqGzTXRj3OpMzJjQ6g/nCZVm/FMs2YvyfcgQK4FjCxgU/oe+4
4I/Xay09DJIYBz+X1QcHknEqTdaN02VeOyO+0qbZ3DlZFM746BdRra3yeTOFWA8D
ZXd0bKvFN3UyO/jcnYnW7oY6/59zlRD0gXCYNQ4LXUKtIaXnj9L464bHRzgg/T9K
P9Tz8/1vRrnVLhdq+VzE5P15kyqnLI+DnQsDNXosQ5sfpw+pEWMK2SAUgCUp2ttz
AbtOeg/zfvBBKHJoCHDsTEBGqsB2J6AwQRN8MvGAMJaYFio1ZxOtGArXc/JJcC+5
UytPPijLPqS+SXX/urieXP87pwpqGr2up6j5ZQQi7X0wzkZQ6h9ffAl4qSJ5ISf1
DI8Lg5ORxPV0CZtfNaG9h1S3qsqko3V5c3Z9R57jTG6Jjv6iUKtn0krjkaVAWFno
oilKbbLbXAuIFvlZ/EgbFIeOApb5auKJVF5vU+ygBXvrSaxn1JAXdSU7xHmY1RYG
09beqT0pAIM+NxecqApLnWShhlIF5Fd1/Q5hF+sKJb+cxr+P7NGhymzEfJ3bnOwY
EemJRtQVP46HU/6Mbka3e21k86Cp6HFwM2Jaq12kFRs96520dfTDecqZUKdZlQEu
S26697Jnn+5LldrcuOxuAmA1wpDZvFUqV/2RMcomdBcHRVJK0BCndioNnyJixLm9
rdFgP2y7x1fE62u29xkIHNR1s86z3kfoOD9SJ11WFPzuWsStiWfn4t8qObM9dXzP
/I9RY/g0FqkGfWToPrRn+uuII1m1LUzQj0Cm6xYCygHb2JgiSZDi144Ob/jctwyE
PLceGpZoNHz64n8nzRP1i5Ed0vYXbVAteV8Wrt9jyY4FmgyVJfo7/KI/0v27p7M3
AomLS1krSCCRDKUtFRXKRyxXm+WTPcSiEcvdQmacAnBBNdTcFE9HlBCW6JWJ6S+J
xjL/aC0Nak4ATS5Vz8vD1nVan0dw/M8dGXLCJS4CMHCLnmbd4pwj3d3nD3WPjgNq
/X4S7xLK75j7hPAfvpdEYzU/eyo/cThMKsaPVASnuOgDQaojASwXCycUIrGZPnbV
D13hlOSQQzXV8ix2cOSYRWCfs6VCOJdXrh9TvVCEDpyqf1ebwUIS0cz2g5GWJqV3
yft638YpGaivZRZX4/IwP+x0jIc3pZec6Scei2wAMsTjmk40fXQqCWeSr3Z90O9P
hpa34tIHrWPdE8EwgpqXhXKLcZenDoj7smnbb3LIiB0ZvSwDCOsAivgKbDXX7yhk
e4YC88zLdHV0nEjj04QdDBAz59WLZWf7nmPCCSyPH0XMHYDPm9Buk7+ccxeXIt2z
hs7pUZS21djKyawgL6PmteH+oit53h+uE+uG8fR/kI4X/kJxg0HCAKCGoVpjBkmw
PdmRRiP6Qsg2GMK/HGBGa+gfzaVpKUyhdjuX2bfUm6IVkIza5ZdGO5NMycyMwOvB
tkgk2P2coOjYGPaLgG7ovo2EgariwOLVSGt8tdIApUVnXMqvLStP2vDegklwZAN+
LyFm39YTvUB0bT6hTjMye+KxKWdTmzT2gBnsihErsJVzH52MuIN6A/iWhzKpwVl5
Xjg6EhQAlPbbgAwZE4aALvO223MaX/bLuhOabpavJXT6Ye91jsKVgnSFKvp5jspT
KdqjDKeoeU1lI9YsQDS9JQZ1AGTF8XupAo2D9HKBo6LZ2jfiq3gyfIJ+MsYUn7gV
YvEn0zj47RXILbkAg8kyNIPAZguYUrLepW/S9n4xh9kJTHm8ijXb6HPwH9T49esc
4yG+r4n9rjTQ1uwCOy6rHp59v5tEVBxghuMg85F50EaKbWiu83u6Svj0RGSS/iaU
xvkAK/FbScVzpDe6dsaU8NyuckCCKcT71gtlwd5HV2uZVnH4C5hwCq5EdfTIpPQw
AJpNgIgm677diS5ySTUFNXImycgq6mzWbh5sCeuikIzPOvofC9DA2nNWmZSXj7K0
er946otvMoEJdW/3joHwNPk5MtqU5LLuyMCcXCSMaH2ucmT4xIh7XSK84WGxJvq0
MG/7knOt0OuUFxDB1pbsuVamI3l9DLB+9e5BYmTeoslwGn3P+QUqbCMK492ZQ3Au
De+0a2GNs1INyKeYz0sLgiAamDL3QgL+jXAW6UKx/9THK72UOniyAgj0RqN9uIe/
t5I7hs8VCA6jOs/0ZqMQWnrY0Fni9lEQlgIhTmhgqjZ6PsyO/Qn+WcP0zTFwevD6
FRhE1bukhD0WNkdFDjk1QADl1U3kIrTfyuGgkzMON3Ga+GDjMF1UcNopHqvdmyFG
wKxR0MCExbrJh6AMrQOY91FIc+jlydIHbGxrYezdLr2CwXmSmdMfrwBUJTuhsEyB
beY/vwehRFg0hVzWmepBCamWSLC//3GZkZUxZcPN2lKmw0n12kjlx/ZIERxBeehC
CW3N8EGqBrTnag64NCJQ97h9KgVP31tK2AU5u6Itiv1e3wciHnlCbF+XseFVTIcR
H/Icz5HdRq7KLfYXvQJArGFn9ZM2ZpckSw/YKt5F/iE1HHTQV7CoRln//VfogibF
WgJYCFVUBm1TGSYUAAeARqMOsF/Vh/ry2XHPYHg5Ew1yGwRZYOcLLrrfH8WS0UjJ
3ARse112GbzbVpGiiSNssJv43NDs64U61lJ4hCZ1W3uLLNQDmvGnvbmXqqHPMpEU
vvETbm15qlnlbFG2HQs91YP+P/N0GbyfaEhAnj4yyF+q6TtalhmKl1LaxSTS2tS3
YqTxmMSlSiGIj8tpCOq/Ll/iO+akxvCcmzetIYKu3cbadveS8lH3wvjIsT5bzn92
b2Xr1cUsusQB+wGR7cvf/rA0bv+p3WKNkc9z7yT+8cpLPJuUmlNLAX3Hs1W1ozR6
2Me7SQaAH8jBXEZjmnK1QCbaQFOJDivJHgIHPmpbRzlMO1+uuJDyuSlYb8BzgmZl
azvNSU9a3R9LlaDfugIuhY9w6tbiO6Yh0ytsE01nLy9gG5Ob9U74Waxk4Xt8GAXA
23pFOSHuM2CS25i87DEcmk9tQ8FegQXa+aZsF6LDs9I+FIDLOyrC5zo/Umzr8LhD
e/7C11naLt/fRpw3vBtLudKPfwQBbX2MyOYRWqjSK3SVp9+sFTGtW0EoCRK7n0FT
k50FpdxablCKhLEW7YY81Ym4bNwoDjNFg6+IZlmaz1uQFCo8n2LVNH2n0EmrQMtf
LSqB+z+GsJQgGcEwOohmE55rKuCc+xlb+dyllU9TeOHcaRu9q/+5R0tDsG35Gz/D
EyLmV9UJCNc8W/Miye/vSUdfCdsSCsVuEKCPCrnpRxCDihy0ONwCc/QnBVvVSEzq
hd/rOAUtPie1E36H1uTrbaXT0gMoH+fH+lp/aE2gGFrlsRyIB4rxtljA/EijdTkg
a6OsUUptetPMxrSzDY+1A2ETt+pmxFqwLkvejSxSG7r93fF6VMAiSBJbchlm3JnE
d0fKHeMZ6Vf2x3+t6A1vzoeBzeeRx9dn574ulFj5r50oeWduYn+sMeVucPHcFN1t
4xQgcxxlJPiZFsrjuhcJzMP78UzQnkJkjFOOxhTuPEgKVi5r2Qh6/n9gYAHVHy7i
IMmGq26BlYFCwwPLcyumwsWzohdUwxvY+RcoRPaaZoouHdFLKvwNgWagFOTjfV+8
rDaMoaeA2vzTH3zrf6Nva+zMFdubNyh7ivrbLcrX345tKq+dNQz3Fj9+p79HcAMy
xT7ORoR96yG0T1/ogN5G115Ze1e43zJNWtJLHKQuWUXb49UfA+CXg2fd0EUVMszd
mb6e5IKgMHzDOsJwbpHcaYdOUtzzjbkeB7HLxJAlpSM6CvtWzVcbWas0dGWgGyJD
Gr5FSdWNsxtyyVX12T/9NtSqOjLlE/AQ4XImlFkU7yM84GAYB/NBEpTrkAHG8orA
4zVe9PnVbcyLFN8egjgCPtAE62fP2MpiJ2YQ0/ONO4oG9IUZ8taJB2FJU1ML5euZ
DXh52Z1O90X58TTpNyolp1Y41W6SNmuVOOBd4i3VQBV+gAaEHDkkwPImgl8d2FVW
Hmzr3PjzjOc99zxDnIgRWBExf4Omj2+UVIeLq8NlTSbDwagwsG3GuBwmwrs+ThXM
O4vC/8FAU9t6PEvtde1LDCdL9kCNq+pxUAYw4/1WK+JhiGu2drhuuWjd5jwGWKjk
68WsG3cnbw68xC6vsZKhgbNK3Wpds/PWZldSlQy8kf4mcB/mD9GsVDiF3A+K6VZM
62Ra27H/beih/5AHwJQNZv69+roUlAEd76TLeUtmjANYhoeI1KHKCU+CJfrvPGGV
O+ABM98YoMTBNNznYj+nriFsPm59P8irHCyaAhcoi6CZG5HPczYEJGlHi4RGANBb
+cCuF2XpCT7QKbrfyGXQu9VbzUGPA/M2yzoEy23agnYKkg6gykKm/yYrSQhLI+SS
h+A5DsFkJZR1/612tXBKwYyfNABFZhamHb/0W9WuOHVltU3tcHv8cydWg37oXe9L
wVvCtf9K4schqlD6kPaAqXqNXlufIsN6irt1vsoKnep9ZNiH+oTNVgyCX02fpmTw
A176iwnmO3O2P8dcRovUilQ8sk6cyqK5go86aGn6c4z4OoO10UKn97sQv6xgZ3Sg
B0F/1/dwqIZ8U4TVOcTi03fYaf3o0qcBzyGYCy1y8oQ1RQhNmAH5J/KmdwSEeD74
1JXJQ7S7MM3xftZHiMD5gIqZShkZq6sOiyIcjA7bAkBlQcdF6pxkn7DVxGplNoMC
yL3okCVyuj3//IMfiTbqJJUq/v+oIZyayx8ymeH7BwYEYZ/Q1aiJAVx8NpYOXkWO
HwSqARXvHjHBsZvKmca0+Bp/RObHXEoMqkcNZcE6xyu1rsbVuVeL2GJC5VdLGmYd
MI14M/bsqxUr+0LE97hFhPp0IDPkHbKJn0ajesNtyFoldLxoVQ6X/cB8X6s1HlAX
rdcKvo79hV2gdrwcs4K7UvfSr47AY/ecsmQAL1gWxwlrBnTmyCwFBUpT6kQ2IwYB
oTFmSCgJB5JhJyR6MLAdBATbRpSuCWYOKwnnOvUZ4/BDW1vnMqBR5r3Jjobay+wh
9UAmHEMf2KhPfd7jytxC89Us1b8Me9lyEAAoaKAh+s11K+6i4gICXHdQi2bhXufC
CEnMPhaT4OAAZCC8Zb2G0lP+syAUuperH/7WvDHDaDAqPiFz+eyIKEguUaXASF3u
p0DBWJwXXuqOvSmidEPxZhp45RtCPxbLbhaoMemMzFPj2HUlemzKm+Ifi4StvuVE
FvnmoQAwWB0r1KaPCO6NvMtuqcvdnbVg99GuVmjH9hxPrAh+oVuUcPIDS9hlTj1w
EIdWaJwXI8iSHPi8aNFGt+Tg/PEbQpIIz+cSTmBANGYTNXSgtmklUpUtiyEjSs0V
HORffTs4ybmtKGzQ8yeRMTPL3iN9xbHR8OwLW/7I5uvkybh2urfFgV+sf43/66R1
RFmVpuFj+TiNojtTWaWnpMcjFbLtYzAVGmagcfKsGaubiMOIj3PoNnGaui7m+DTa
thpP/xy4XXOz2T11/dS9U60QX3cSn/v0eQYUPakd9PQP/RiyF/8P5zA5MEQA0qd1
rQ2o3vYRDAegoF9TA2qnettybYXgHHuPTciLfDHmKIF/b8Mh6w3da/flXjB5LPVn
wxrXDBRvEPTH/e3aHe39OddcaaxED7lDjzBh0rGR2Y5sYFByBYIFeMCLHCFV0wW8
PRd++UTUB9hDMLq7UXUrsGa0LDj8Fqa4lgEq7KAeJ679zzjh2Z7pNFtPby0qFU5c
PLXgRfWydhZqDj8oYYKVEQo2EIKjybvEFPdLCmWebHVqQKJfDDzDh2aOqwA4ukJM
+k/9XHDLywRTs/jialx5tNVV93d7cUWwULlY6xI/k0WtNz5KcD82AF42JzHMqNuw
FSeUd5XWkaODMePtan2/LuwFqeXRDIp7xMcj8sFrJ7wDfbK4ulDz3r4KqZHJlqSX
Whf5i2XeoXYorNlyV32sdLABMasSpPyELqtlLj8GA60xcwwamB0zLwwFpvCeK/Qm
pvJGRR7S5FPxXspESvmlzoBG1vy6swNtluDM/cgJ4V0Z21id3meeYxqSjMFaJxfb
1ae0PWaWxJ2BWGKEwD9NND4oZK6VJIUw2YSoRO4B4xNos8k2PYNs5WMZhQnEONRg
6YRqV2v5Ccr+6YJJ86NlLxDTNHRgsB0m3XLPCVYG67HlinEpJK6HRkB99wGk0l1i
z12OPPQHLlzI/lpe6NFeDCsVZoRkA7rRFo4nRxJEtxnA3IWaQ4jd2b5LnFV7fEE0
8ylWgrqBPE1okDSoc/aUep5jcWKagalMCKJpR4EXnlQ5PbOruFBlEeqCxhZcDFOY
//UGXGgigo2iEjJOTvhkiQZVXDcTaxdLdvJAKwsjgUR7aJrB0waaZt3bnt+Ag9ce
lBb0makslo9zNPexbfD6ZuJ+RrMLrzNjy+PwHAvccpH88/e8cXE2urhE92LtWzcP
SEgZcttxqF40TT7u3/ObMBLzGJCIWNDuMuiuU9mgKiv0XbZoE1jlFT2IiEiKV6F0
DTvWEfSCXVhtU6Kl94mHMVeLKaKyWt1n+HPkBXv+jb+xa1csHvFI6uu6RTF/wthG
+L3dkz2O25bbJwV1xFAnnfT2OJPgsHeEHJ00grKTYxPlMAalylhVJxINDcsNYjoc
fyfCviX+Hj6TArPLRChMDw1MFKx4LEHB3rczQwxt+XMoSSEgoNMGHgJTl9iDhtj7
4k70iTdYfZajAvxXcXogDA85lzTr5W4tRPxk3nCQcLwsZupxmvEYQMevMxM83/rH
44WMqcth41haSPOXD2V2Pp8y+ERpvcLA8UlARq9p+bF2QZvENr4VBkPdpQPSSQRu
HNmhKo9GjtM8pZ4slUn8epkC0IBZ9MT/1ui/sTClEw9CWuRJOdPBypqTiPKEVSGk
+nNifohqUINdrBYhXDTiCsiQmE+K0BEIeVstspklPGg62xj+GszKYJ+Cy72QRNr7
qspG4QWHLIRdmj11kbFg+3E5xB/PbnQUWuewLDeWgjRgUbRL4Stzz7xpY/ZRCZRM
nOHceJI+f/YnTvVOi7A3z+UzwPW1b339avGgLD6x7bejp1YEBvhrYwjExdOcvlxO
dDDWsV6nBWL5oQJl/JxF257WltBDp5COhUgwq/Pvx85L46MES7vlfziLSQF4nk8R
5nQa7qVS/skOngo1y0On3pkYHvhKU+ZUh6aNRanCDmKuO/pJNMYZ++Kdo6lQjYuX
OoL7P5eBBNl0l1IoRQNv5Q5mT4hmx2nnvayvY9jruXzSHVN7hivXCV64WmHKnshV
CbS82gSi9Z9DGRpy4nL063krJTBu7oW6u1JAm9ZWvN/Ru71JVuIXPpOAGk9GC7th
JteXA2LBz3jCECdreFBAkV9NzOXn3f4wyJfGffwUqSfzUnt2xGsr28QpkUJlhfSG
zTINuaS6/o4NxbTonb5eYPHqDthJZgQnPA5DVur8Q1kNaUiXpSC/iabq7mp5gyPp
lj5Y9b7Gbfm38FSAEQcZfVDne5jsJQWYZtIP/hfoClHhglm8ans/+vGj9nUdsf4U
6YrWo5hCkhKBR7vLpAs2WzuH9zKig6bCfpLSMkOOCwdcAx9DJEUcnviwVnKjfiE1
mh12j8kDKhxmU4Q360BygoDhPAzIrDDC5WkI24nfmpDkdcyhy4iRJ3mwfe3uF+pQ
ogHt+9rt+DXREio96QwTDq4inhIl3jI+4E8cNJ85zO9fvd3woZgyRGnIrTP319aM
NfR8yUavkOXehtq2f2MDWcif4Iv7BUp8zeEB5zjEFsCH5eaKqdGTIT5/qNhp3750
ZdGdrr6thF/mu6gS8efUrzHUf5359oAVyGg/aUj77X7Fx7cUbtqpBKNbYgZAfq/7
EuNoOmz0Rd+xlonFq3zpOvqNMNxEI/U7EY/qEU1OUh2VY3IXlmdzWKojgJPg8gYe
Png+kQLGU0qKMA3Avb16bbvXz9+DDwGQsveSHNC6yklw56fZ7hqiGmbqAEeY8QJ0
SPuEsqwbXhpuT3kpljmA4zKZ8yo1DALnF5QKh9UYWn0lTfmG4S0lm8Il6KDblxoY
4QjRUKLCh7A+HxTmRaFcQllEFdI+Woxm52qO5SvTmcf2qeF4fjeZd44/dDdm7Ptx
O364c/7pS1Og6jETo+6Cfqs553QXTyBV/UhYof7LnHWdHSrEbowW/02Y1mgmLh5U
CeSZBIB8ZCjRdWOyQ1dOH2KtKhrmp8LwGthG+iod9GhMwnIgbIGoYFcf3mkHh6ZG
4Yza+09qsEbxTIBy3ZGz92HBVVyOtbJVqfD7qerGVzjf/G9+qE4r765+Hi9Nccr+
BPu4289RqSAXv37PRn+GxggvjLbbyxSmUq/Rqd/onPKH5f3ftazP8ygaf9mt6WCU
lWg5/vnfoJjMkEVNX71EswTRY3HIRoLqculZKg/nbhZ9RvE1k/uG7urKXzkKVXeV
x9YifMNfD24QOSE7unimT9xUNk4IPBmXKPwREz/Iqfi+xsZzdWYGTUfKGQjLtSZe
d/KaYT4uv0swDVn8SkokdBaUusv6Kj2ekXdowinjwmIcgC5XGm3vLvQC7flvVmks
FbrXK8lm+Znwmm/1H8Y103ZGth3EJKCpp45+Uukpk4F6S0TZ/oQrXY85BnpaeKS6
pHOMyl78399HwIPRfuk0P3SVm+fXsmPPL0u8JQHXvzg5muiuEZ8ydcS5DqWTqUsn
odngbrOGFeuhzjo1lCTXyRLdh8E/egeJ/7j6WyNgctsRDvBqb1jP0Zyd0mb9eHns
LtNVgWwUNiAXiSB0RF0meU5foGFqyqS0FHiOB/86CFhOXEbgK5z97d4K9ZqNSCLv
nONUvSRE9VjWoGPU6vLAtlhwc+qNho2n2P70nAf4UlHFhF2bUOQ8MnIeVUlnD1zP
U4zwzIc2LrVp1J7adhv8R7FkpB3EOJjIG3+mDUvG7S9dYlnAoQyVk6oHeog6MRX8
PQLp2zr8jQYoCisa2+X6Rv/6wSEn3RBix4ausvKG0M/93pto0yAd/T2apFC9+a4p
1BWi44CTiuP30acSRuKn/ZqW3DGMboAaHeSUh3BqKfotz6Pqoue/SbkC7mFBOqo0
P8Fwea1O77IHAN5eZEx/kltSDzPxKAcxAvWNxP41p+bZAR+7AZ/rhCF4dtKA8CNQ
sNNlPP6OcxmDz9unvWYqIrrICyB5VY9K+AbK5V7xtM0xAnBZK2NjTSw5WXB4mjNc
ghJPVF9tzt/LVFbxqYae0fEHDAFryooW8n5CstkrMw1v5Wss50VIwPQDiZCKpAxw
Grg6EWkRS12af+vlKc+JzZ319JE0YELSSrm1T1ut2njITHYknD7VUv8PsfahIB/+
xNsrCxCYhGsMy7O3Cy6wmTgKiUcpnumWx0v6qfDMgLdA93xxKk5xSPukgaNdw2pc
suEXshfucOxCknaSn0VF1VwYxUFedOWxQyPYtWBRv5bCSn3DB5feqsvTGGqrxJoZ
6QU6+siMAYlLCjyrYOSbXtymaahro90iAPhV9p04APDscLWTHzxwc/pPzEKN3fzl
7I6Uy1vSVKtEH4GrMHvmwyjCyILzC/5XxF577UVc831UDlz+MXg4uNXeZhfzAbQf
BBraGzWI8p3SRysxgGqDtSF6wn8PoDLPpP5hWXTXAVRHsenNpTYRJe+Kd10/kx1O
90+Sia/+Z+YOAwuCcB2MSNWN8Ez2EvwxYzk4AQhm5JwZdWoyBT6/Nf83vFgqW6I/
v4EuGtStfDQR5BjJWzQNZwkWa4XE0il+x1xoEOgIFHk+HV13xcWIsR/+2bVoFJgi
uZZjQO8RtQn3rZFHL2v7q+gU49IgZKkD/Ao7Aa73EtMWAP/SP4inYq1HFxsTKokq
pxSXx/M8clZTRVG7oR+iu5zzqJhxQ99d2TmucfCxQHm8aebchRQd0TDNMQi1deP1
EPgrbcpYqxhTuwSLdCbCJObugInjr5lc36+AJ0JMr6WQD4uEtXnIWfvRpgHfb/tM
1e7+NYiQotRnE5c/Xjla8n+Dyhb7GPKWUpm4zflw3atTMN++FyCsg+tXFTOTZLnN
fl+is5unhSWw3BKS+y+xTuHjhmMqKfVAYH+wn+YgKZRRFuGSHJfLO31V0hunBAIy
x1cblKIeYhtUsBb5DHG/SiHtNb905gv20vHP07U0WoM2NaNoJuB0QbZJ9T5BmkbK
hk+Rd4akdV/IZufeoprTlBUsBMTlpCzEA2da0nNuA4BCf5Td2iLjEKIiVCK1CvQn
Lq5qbv56YN0E6vepM9HXI+x8vDcXsTIsoeSghvu5OyY/n6RYeimFeoPIVj/iSzjc
KRTTc9fa7Thm/CXfB1VkYZQx3M22tqWvPJ3VJ58WWJo7mk6C2FH95D6x9qSlggdA
1tDSgKD5l8h4D4d0KxARW5PFm9gsTLHZKN0PaEEtIQ1Ax0TU1avHKMfM9k46DFV5
ggScsnK9LgeaUmESh3pMtDCll7y2ExUcxjG6AaAdm8+AwFi2OmcjhCb3Nbp6p+JM
iYwFVgVS//b9osOPIHU939BvBFHqlU1Y527mbUvWy+zyH1RW5KaOzIdtVk/puYV8
LRWG9N6m2jNPVjsgLUpB0u7p/jCuFsvR96skogRZuiAXPJsr07orkXEIGT1eJ2k2
/fbxUQJH/geBUUsPqQQG8YHHJdqSs39kt7TS4lhc+VPdf5bb0YKxvMDUiICiTNvh
JErSJSpTwPrzCrW0PR6vTM8jUEttxm/xS5ROdXkDiHEBXJuOpAsy+TaRriA5Ox7w
fiR5c/UfKLzTLM0xxSxxezswR7p14D1zYzmSETgfhDeeAzss7FpsICrci2yOui0m
0pl8S0KTRjOEQaDjfgiZ2TTTZET4g67uwjsEVB1D/x5D/k9Bd9SPXDdQou+Zn8PL
QK4nAcy5rrXmzeLGMoNyZxOC63GJ3d1uaObrjH/0/0+1t5bN6jKSrUY1qrwirrB1
dnLArt9wmglS/ca5inHuHK8e/WfieG/NaNL8kuPdnC7B+X1KPEZDcjDFCUGMzIci
UZ68/eOzDs/zXW3/VSCpFX/5Ra8FB+fF76u3ZBI/SJHK+CvilBqJPSBpWznrJMt9
cuFu3eLHlFiRPEVj4jYx1ftWClFm9XDQA4Q0KexMahPi2juzlxcM6CF19tO5V1HP
PycuHUNKa9KUNRBSgit0MINQqOP7EroSuM+PUrZVXRgYtU1DJ+TLAK3M29Z78fSx
4BF/LowD7eGg+xopYa+5Z/5A16ZbrfH5SdZhLnmNnIIpDsBySPArx+uwWZkCaQQ9
HaQXXrE0UmEldBjulRNB6MqIYlVhXxaAhcwh62kBtGflMryfZlWPP9DFr6urtj3+
9bbx1fjom2cVaE3eU9dAcEwn345zwrM8ztDxuZNxC/WyvFGfk+zkwUU65jrjBIgT
p4BOdzR+VUem6igltFhJ6B7WjthawdF6Sd+wea+VGeYgUtphVOe27AyyRySpmP07
u2GxixKTSiMO7pwTYeF4V5JGYRevaQMiSoEr9dIkHw7ALViObStdFHbgvmlWfTb2
hX2kqL9Xa98nGEOhjuvaP5K2xv/tReq7s6S7jR4P/XwgVgav0mvcgL0C/O6aElrC
QIYD64ubIp+sBzt2xnySTg1EjyMcTxKNUi00WNhFUianQYUbo0b28RHPSnPYyoQK
4M4BrNGbuJfG8JyyfzrvJFiKunWuwD4GXHd5AFhY7bpJRbR4NOLgqtJzpls3bazL
UpmKWxWGbZU93d2FR1qeP0G+f89F+t+hopMBXYsnJHfhK3HzPdojmU+Spo7Ik4//
2lR9uTkotuzRfgimt8Nwu2Ggryyk+c2LtLiPqIbUcEcSGpBe/iCOv3fYH1N1DhbK
JUjF2XFK1hQUcig+teHiyquRoLx/TeXa5AQfThcDksAvD2LG0lZR2SI9R2nJ2pIP
VXur9sCBj7Ju8ok9xrOYUJG04YqFuYY0whreOWtIgL2Z8uii5GKbb0+4h7espHGQ
UvqzkuNQo9XYVcIt7vvpbXnhBEmsfDxApfv0Jhh+iX1WfjOF3ZjMJklbIcNSsW8Q
T83tBPDTGQqFMIhXXGF62WL8EpcC4hmpQ3qPCElpknhcf5dafIvhm8e+rcF4AdiY
j2lvUBR/6MOyUVAC78gX9tVczuq7IxAU2TgyIV+iSV1wNjSMhbsbE+5korfyO5jo
Ww0KIA0pHcVymQVRmkr76VxtffS41CjHvX8FJ+cGx/TGLsQfWKes1OvexYsvfmgK
a2Qr/ffyLsu4kuTSV+vxvyS307QdmpGIZf6YPB+oItTD2jyYXNGMzbCnPtrwzOUs
OdX9w6XrQnAOT4f047jri8N/Yu+XKzKni2G5aGwvLx0D8raHG+3NiMzpFf66aStP
Ooe6dDMKEROikd+jaZYLoF0wJkzep5+k0uMcd5h4tNT8CWMaBk55iN768r80cHW0
4QK7l/UsMT+/r62+AICICkA3gwx47vsLiPu/LgOaVvEgF0iRtzb30bLjZBrciVtS
aC7g/ykiUg4ajYCeGOC624K/BKUhzEPc4kiZBa133wpDsm24qRR4dAZGCPW4SbaP
/iMYWvpQqi5P1LDmVpOSHtFW9sNjNs2r4gl77g+8RlSGuvpn+NengUpRUTXE8Wmb
kIFqXdoh2Pe9Xu53UTiclNXY1A2wjpY/DweCOcNqvMsFeZcg1xWtpFe1e2m5EL45
eixXvO5TTYZQI43uDjW7LvKjWADQj33QHexqJ+v5V9PnHigJUEN2iJRCZOLAmbPj
ochi33eYIfCZVt/MBdi2N4E8vVfAmcLib8KYnwacn0e44rOxngeyxtDXyNxL4O2V
r6OPPgXF2ZvUGFh0I6lyFI42sMhNvXg3V8a+DFBkYEeGn97S/Mrfcs6BQJwxPXis
+hBhYSZANBwtOs9KhXJzN7Hp3ZymIUpccfG9yzqrnEgFAdabpkZdFydQ4o9eGIa1
0dSYKBRBVdZww42+VrW/t/vpYD0NladdfSt98aqtB3/p7dNpmwaJk7rMi8dhlUX8
3DkR5b/FZmch8V3d5KyEqEFHJ4QJiHUZ+V2zTX/93XLFi69NQQskz/0PH2wd26D/
MGnxSQC8kzq8ZBwjcskG+Ub3vmSxAXHlI8DlX8G6ptJ4tAJ64NpD21kuk6dXYmhx
LcoVehRHh7RLlUaxnZhYal5FsXTUnn0cxWrVi90Ouk57XP5XzuuakUPTc3wg1KmY
jIZF32nbbx/kRhP/7iBIsnu+QqNO0ufgUBKoSTdzt0cubVuOAR738CKpFW6YU5mi
c1y8n2kT51YaF1oOLFNLAD3RFwa6iTaDK0E032bPszfpiHDLWUGy+TiZkeIw5n5H
zM6WdSP1t28snTRJf0QzAr3uZX6ajxQ0diKmzYmuH8v87MAzQVj2GqwuirOHCPFu
+kJ3ND7A81LWCj5k+Y5+JP7bNaBevlnlJnTHn37+0tz9fW+5I3GUlLADYbQ5Wc5u
GTsUKRuWbfgdzKs4jsYPpb1vJ+yQer+CvJuWSfXu/HJ5g/4AGR+GP3nCrgeqBrls
nN08xMY5d54ouEb1DmS475jboGtTr4goGRwB1Iuvzy3MsxM9UkIF9hfgCtXsiirz
VijOqmdFi9qAS2Xk5bomdefo4pZNHPzUTZ9z3mY/+GWHUz2xnH+e9O87bGgonAuP
dGrS/VTn+zuhT37L8O7GBs9iV13MwIZGm+zimYH7ir5dhPWHD5zJTsd8YYnKIVi9
Z+dGuTNwc3pbqf9g+8JmZXOFud1VVtbG53mxTs8YneVbKXOYR6A2IODm4iL0GaJM
b73DD971+oGv93k5Hwsmv3twRvVUcFEQBTI7y2uRnaYX/gDXFSVYhMWRakpp5p7F
ceFdyFVj/aQz2A4q+ZekVBl2c/MY45F9vt6EIXY36YuwIJcgwSIR+EJqNaf/N6HN
E/felcrmiodUCOU9ZJe4zAJltZIouhrZVD/wlCJ+vbA3J/0y+P8+xtl0Bcp0mUtx
PCHysp+vIfY0jsSpFMaqouAZYh4q5C6fp3xQqyepYNQjkK16TBvuyMoEjr+edh/4
LUVBbIAyw2xBBAsYouG9zj6bLVufQQuqiqBNztY0MT9v+b1f1JgwCr/KbqmazOcY
VP/c0G3GjxZo4PvZrsPI7g22UAcPaMfImTJD+Mgh+gHlPPcye6gjv0PiVAvP+fEG
jzz3r4cCuyhRs4c3ZGwRrt7m6d9nQ7O9h0IxyxoqJiNf/gCdugMJ3Q1wKH/sVM56
kanAcOCGk+HCBU0DLlL9PDaPmTI1SOTRzZ/2Sfa3VBqOcvotiPlY8jKin6Y7y+Qw
I9C+lRxx5A1fkiOkMVFwkVHSu+8ySqXEIWFo3Tgxxdh2f26XoPawjMyt1Yk+b3Yv
px2v8LAL+kjN16zRLnKvMaA+ZPAfO4lMrGraXrDn+VoGgrrTcUriDlz1LV3J7sHV
VWh1n7BuTcEOMYjwLXRV5uBssTfOpT7XntV9oVajXMFiAa1B+f9kM5nJekWVRCAX
52YPU5OGfrMfV/QOd/Fu4qCArtQsofo3OpRwYm64L65Dle/dZE089kGnCwfcj5K6
AbrnY+P7VidOwR+Ph3GQ6f1/q7OVuBSn3188KsmgUAYRO/2JEfAd53/5MHWbelDy
l4HeFFhQ9oF2MCP+SUlBDpK3i/rQOXKXJm2IIiBOi6boSQwbX6jddKZtP4VlVjfC
mkkWVVgUQ7qP2xoMYSenAvr7ksgiRr2M9ckxioFv/0C93Tp/OSrY3nz1+P1fEZnV
9D0FY/JKqgyPwdRA59jD5cg7XQE9wjT5oCjzj+2CkOFeM7x9DpOVIl2CnqPkL80R
WoQICqYXyAF5kX5/gHyoFIqQfTwzo8Ivh2mnvh363wysmmpsHtrFhp8+lDwB073b
h0M2YNwikSOoa6AOA9FCRCCLTadzrooG2rEAGXQ+Z79srt/mRWpclqYqJxGC8a3P
fR0VAYKrHzLxKo23RsEI+OVW50jD/dfm6QdoBFmV1GyFqCu3gwdW6AmYZuoWJnW+
2lrfk9mypXVBZxDsEOtRqoVdesbiaT5KT6q2S7cZaluXbIZVtSiL/CZSHz+1kfAy
qPKUkE9WLuSlr4JuXs6CCkioGOefD9f8/lT8RhvI0APo4HdoPCIuqv0a2RsUaW2B
b1nbVBaEkzotT4gj9BEtJ+kHn3FFZwuMkr8IV9pmQ6nA6baDZ/2tQQUlOqHrxgPH
RdBsI5cnLnc8XpSM/zQHg4uJbWQBrqwhJeSK3MDzXV6MypcKp/IW5ln+HUCDPqSe
qSUQvNDyGdY1D7aA4+Ij6oCqtP9FIegotmo3QmHkxzUhZ4sU4e2kwZmYVM0FU9me
q1kQIypsa8meRSEZ7qDU8HXA6AAWISboBuVgRGppmMAUJpE1ej1WGoOeAIsJ6YBk
WewqoLXmRPmNeqmYpzcAImIbOFUtKnLK2UfVp6WEokUsueTvpblbrM8O0a1iWMvQ
cVim14qDcbQ9Wi7AWpg0wlKYUxhy8mFkx7rUm+iezAqxCwU0FSa4GADjspLFcmxH
DzGwsUVaGFwk1eS4rtFWNLClnlzRR9DANQZunzq4QoUkaoR6zYd3xsGZfYjsbWg4
64xfPR0waCsanK6NYSVfOqa8Qws9LEiSCaB6kH0HswEVf5anXHDQ9a+gOeoDcfyH
uEw11xjyyn9a9DX4I7JbSBky96uVSuCtQtM1zkJ0qrgI1CpEGjFGMURETqi0P1eb
P86ojniZgJMvhQ3+gFislDv2rw5gd3SNn8OL1nvnG32548jDDVkCyOWtKoE/QUa1
i5ruoMAJD7ApCHePe2r5ECgCRkbfaFOy/QtZaFIdLTZvs3hGUn6rvW05Sf2mrfdj
67HwUZKahDOdK7UlMBgPph+S1ijQcKrqMQPElhiKCUiu+evJvyVW/3AdIo5cbSfW
938rKtU360Kc6Qviuix8H0A/Z7/IJCY1WL9xpouBIbyHegcKB+/wIxURq5/1E84c
sdaLLU8f2SOkufHjRuxZ9A9DzEKDQjT5WeXIfs90OnOet41HUWxeSR+/PqqpTuFV
l2k9vxb5VQ2TsLV0XrX8iHBzuYuecolyonZ0/GaTE/azn3sRZ4etRUahu+INF4Wh
Hqxz+j9YN86JDiD92frtmzAfMMw1T1ot8/I41tDpsZpI1QJBPymUgyA7K4tjsIXT
3jo5el2f+/AH1bZ8+dh8C/KpWTD1vDiq+Pj7giWEy7ACCKKoiSvmw5mrwcM7ohxn
EE9QE91Ncad7iBLif0d7ecvQVfd347RITmkk9HXT8GgK+4E1Q5me89VRg0f2wdew
lsbGbBXXIJ3vWfUoyrL71WTef8hkVaio1nfIHV08bMxCcY78s4t+rcoB2Tgf1vJ/
1SHmGnjoWGDETlWrKhmDADylLNKkX+bqA25q+hlAc526OQ0OfYolbMA+fjYSYBzI
avbYw3sli2lZG/iDaKoEh/obaX92IRkirbCIxBBsgfyYROrfj8DmSJ+AW39Pkm/j
Y9WpEhV0RcpL2njOEOMkfXnHZQNhsfW5KeEDTbOgf85oY2GG63Yaov0MFkyAZDnG
ESU+y2JNxYsEed1OCNoVDZYQ4qBEDjshx8WZucPSRO9HTnm68tzymOnrs7lhsBGf
vK419eWS7EVUiWA0vedHSOAyUJ4G7G+NVJRZZMytg7HE6NFwI/qEr32J3Psft8rT
T5l6D9gMb8dyN6BrmAphi73l+OMo2YluSsvSDnGYOouV1DntzvaA5ILtbYN1bPAy
/fwKml8sldQQlf6USeIhKwfRkO81TqD2zfZBa67aZ6waYy2NHDVr9inztWmDdwUe
zYHvuY6IpSmNZzqkCmEZUT7f2oYetJBIXpayA/xbiVUqDrdb+ZVWK7ND2V0Fz8x4
bTE4t5+SwzaeiGGyj/Uge6Z9/vov/3wCF6Hf0NzT01BNnyJ+NiVsQ3NXmmr4oNic
myizIbEAEeCds2DAQUwt8bgeYln5wZP6auRGLCMsxA4fQ8NECev6Tk9nti3rZqqD
MwAunLp8wShU8ft1/+VykadcBNLjpKgKXqX5jasLyDfpNnN1lr6UrcbncPM8qw9Q
oZ/tOGTKx/CIaxqvPQJb17FfjjbvrxxLB6Zvq31k6OEgSe7K+uSwHINevH6m7ovh
HDMDft35uhCy+W0jIE87ff7dhCrCqSrcnFq+LoLe10jwu3efVX7xM4+vUX1Do6yc
M/qjHgs0SWabR4uZRBKV8KVGig+GVQJWynNayc4MONU+MFtcFHVbgmz5eF+WnU8i
DZkrv68iHBfFfsYvSAD3H7HEGw40oq15Lp2dJZjM5s7Dn+2qU+LvJ3asFX93Sjme
wSrPYkwK2UDg8yVlchFp6/SyoP6zUh5LhB6Dc/bRV5tcN8NGThqXrURGTuOMyXRG
LXHhhEhMhzBqKl8Ljh2Cu46DwXMbX9RgbKS8KFAFxzKPluFlo8nW2+OjWi/wYtCp
zira5c95TkkbHKBBVA3l6+AAQqaUGMUZ/ke6WmIcn4v36gnp1L5VX9XVGDV1dn0m
tYuWXDf+J6L9DceB05gXdviTLB//b0wVI4A0u3BqLcJD/H7awAwfPuVYjbmmbTG6
Mmj7JgfqzS452qBLnNquB+e2hexx1vIIs4rrzcdlmswUvE2vWfLfnpW3ctJZgUAA
2O7k5/dSa0itlwbaoklbgDMnimCg5PNgsiQbKXShcLo4kutnRmVONYx+3xIMaK8q
fKlLM9v40NL7fg67Qn4zOcc7yN76pJlK/QrvMXvziTgCb6mmjhBl9H6wVwLMUxCc
+/RaP9o6pJFY6tyce83wYE4JsOOFWHZIObcJ00vm3R0Llp5YSSCuunxfqK6sGLDZ
6mcSZY6NLYL21fdykani1Rd8cEAYnNAAPexJfoNVwvTspMQlpyI42133pKZVf/bC
2ChfbTRjkQ83q/2WRpe3Uv64WG+amjJf3yFAD0ee8UgaSDIEfcsX2HeB7VnRSQAC
xDPnPz/p8Ua1o6GK8RPi20ZmTvi9pu5nSrxci7XsEEgIIFH+cVm/KHx3l8j5KoZw
F0DgbbqgyKlki6QBE535E2SDUydYM5UPgsKGzERCyQanJ90L3f27on55/FVcrUKC
CEJUsKyBaQxGhh+2V7uhdFHjBjRmDHVL4J7tqv8MUQiRwJbuR6P2mTtrrYqOEnc1
Ah0zriiR8QfNbxXTOMzQpQ8FlHlrKRYg1kWkzKh2qpnOvLKCva3AhQQCnsSqlPyU
MKrVcrO2O6deVSwNwsFdijs7ZX8Oo0EShDmDSMjdiZu8woiOhP2LfgcfQbe0kLdU
pBU/G9Fpp85+H7RGAZbolzF19Az/BJBhfYN7NS46Y6vpU14arRgP/Ha+Wj8xruOy
rjt8ey2p0qYwEwIWVJWM4dDfxd6fOn1YIPtlMUDD9uaYUOBnVnZi2gZfEHjYzL9q
NEhtNlMROr3J11f3CgjYXctw9q2mAngReeJXYh6df4zkGkwd2A4vMlM7mFS+EN/g
N1anM80axADQbYdIxy+7CzF/vDhbNoDfPNn49ua2yUQi17pyR2x+mqYPveP3uLdn
0/5yojr5imTFkVHN7JypXM28WTkHD542LR1qXIr/nUdCezPHDBMKggVomoYbuaMO
O25pXoZwGX8qFcMEURZFkBs9ml+XzcAHUgy9Gw6vEAk7o8rJYOJSpNbNEnBTAany
PwR6uWSL/hRxmtLjAcENRV7dHn+K+hDIaA5J2Rdplhnv3ihVUJoXCTrGMOmnAHVz
S6QS6Gtii300CWrNragqmeQnO71VW7bxVNM3OdbBxLAysMPYm0tYGC4FcoQuWg6d
mVnZUfzGqCQMBfNtj1pwd43Z0C5hwF4d9gk8lGSEkzSIxtYGpqvLsbxWpEHYuhjx
KShSa17Jcdb3ZaHdQt8Y0TNz+6flhgM4oK7GAzbyzF9KgO8JHSFFn388uIFB+bN1
3Tv/grg+9+6Xld3qUR+RgPb9Qi5Qa8Ha09UF8ynJ2/TeJDQF4kIVmu7b6ps0530i
I2ZTAvZdNwxasihuWIVANMWEG620ct4QkbeFIA0luxtaTKNxMPjr4WllmTlWIgkc
ThkifGrFscGCiSyRy8T6mvJZdsB2Z+kCIVJutjuRSKWYLvPAmoVjbuWFg6kErkwy
6ya7QbYyPTPgNrsSGwMRsAqLnNLLeuolZpm0xZJBpAjM30k0tvN+hGKoRhu4WI/h
JL02Rg+hsFp4eHlI9yn9Z/NCH4/RSNGe6ZC1xUKEHTTQzAzQVQADBJeSasXyBRok
aDomr8UdBHNP+RV8oOkjE1ROUEQlI2vWU2SETVxLV8c7am6g39M6cX1I4iCDs77I
0AnImWzfFfmJ/H7q9QF1NilI2yp8cs1UoVGzP05hxgm4nHEcJ8HLmGEea3aUWiuz
dn6Qp4YhfhaLnauFqzwRsPhaWxxixHJYAyNRwERnUyBF7tRI3YUCagatOEzK/+ac
gQ0L1tgkZO7r5t2BV9h7W0/uda5Ledt3QEHI0BvySS7QrsB8nvB5lMCb1hIbB7ZY
8/KGmKFcZqwI6BBXwwR9q0cJAjpfo9Dwksfd8FbkAbjmXKHaRr2QFFX86xWFg41o
6rB3Oxk+3VMyvw2u0ev3f07YP2td41tRljIYzqKUY85nef7xP9KQ5W2dMtHrWsfk
VMK4k7VA+pGGYa4ZIRMttAWGQh/o28kjn1GWq1pampRoQ6YleVWJhKDHbmMccqK2
t52wA9j/hA6a0BbG4PGhf3Wystl/3UE7h7Y8uqRTx4J5FDfq02EjKtJwx5kFG5z2
TMMjd2YnIis/35ltj1S0BZFwdtbxIYJo2OiXSt7Bkaq/H3Rm8ZPEgIauIU8oF5An
bTeR0dm4cKbZGDigZLnTf6aCLoSFtP6kexhp6HXemyVehbtQBwATjyngMDqwPdje
iQ7m/8vC0K+Q4NsZkHedGX5C/SJK2shCFXs5wFap6KQhk9qiaLNlWdi2/5k4/ftx
ucbZgYVo/wPI81+XQhOCxcY8KNBAm2QovaP2Hd7DiSSdOHyn0k9y1n8q7W5kBQwF
h/a63fgH/Ly0H/HFQgcTD8dOixfuFm5Yym6U5a/xx8X2W3lX6A/9NtTgBB2B2l6X
GItQC7bk9I4cCLC1htHI9LM9eJmjkB9nVrDf6BopZjU5PKc9mkCQpdJHNhoXPyM2
k3NXh3EzeUS/7q3uxJSTTgpnVc4ZDP9KYbbqkt+A7WWrOz0wGyYwdOT6DW+jCh4a
7dRVpqyCYMFLjI41zHiKUwPmgE1DVpTS4iZ6fK67BXefNIdNSs13RP4P6kot6i9G
kpU1oXe2nnJa3UlMZHMQ2uToIEJu3BvrSD2lPboWgXUuguV856OrnI9bApnQe6Zy
Gp/AeBH6v+7HhUi6k85hNPW8gpN6cVOOV6BQGje/g9PlgAeNGYWWJ25VjgMu+qDf
lf0JumN+/YOccK6hKiAUGDr0MrIKS+0NIzrdS88KgVLPSiROFLBs6KrhtYhL4ARf
kGpd4HY4iqh2CBiYReBVcsCqro/0RNyEG+6GDk8lx0VQA4+QuPf58axHEHKOdrQR
SBMyov+0r1CkA7YvPkbcDK2wzA+3j8/s6HiJoN9qIBHBupRDZpnDQtr6iHscLOkb
XA0yvNmKTOucvdTIMYQknA0SRXbTpbXeBvseqA96JRkUZnhCKHTSuttg63pKvQKP
FEaztBPTXjWhCTJd3uwf/nTvlL+pi7Eu1o40PcDZWAv5JpxgvVcLFzUY1nl6vS7a
2kHEmvpPE1rW6ByzaLpwCK7Qo9i0Fe8wDIP1rXKcwlYvKbFXaN6zQLoC5/pnZSvH
4gWaTc2YdeGs6S9IrYuyHk30BSzPR2qOHemXFpLHfV8IPz0Oml71QvmOpFcyCPg7
QpC4ZMKjpBt87zZmkhec1vgXtGk5DjhKqvPfSFk8d3Ensxcqn7tKygW2eXk4z9u9
RI96PDZbZkoZxQmlqBW+1lwtLhEO1pq8ar0TaHbWqb52b6abK3Ob4t1ntwkmN9MK
dz989VQD75qgvvLhILRmEXNwRhODQBCUd8x20oqokMus2LddQ1gju6wArSfB82ur
MJHWAVkVy2FFGwGrILR4fkTpKojEObTd9SeYncqAAmZVJtKxyUtn/vB77I6sBvHg
GiOTqqOBOhVSiKl7AhvYN6kSrVXbXr1cchugKIbxIndkdjjw6XsOi58uYEHCFJ92
CsjAla1ICccT1513puTcPlgUMeHf9By30TCiJgQVULXEHOnkeYcj36km8p8JSqej
AO0uRyaO8r1vXjT2b7TZUN1vgvWo70JmJYSmiAJRw8hbRuavfqlk0ciA6r4JeO5p
1MDW9oe9t3h2K9MCIRd3PWs1+ywAFGiq3y0LeKLIa3AU+kOO+fnSKpvm0snb2p5f
4UquuGW0WuNEewamD/VHG/mZ+q3l07I2mSkN54bq5cuhOTTkptQiCxUzN+BEN/Dh
8cXylllkAGTC/1AlY44wYnaIRWve3RchoGKSZiQM7gRBXXZ01Cr4+T5U4HMNl3eT
fzk0LSk0xWFk/BqBEGz/ZmGgDHKWZF/X6X4gMZKY8f+mowIzuijkznKmr/xGU0Po
fn0V7IdKm2sU5QPaL83YsQQbuQtASmo3xuK7t5jGBHH48T3B1LkuTgGCHeHAHlRb
PT/1+rRWblm5dgiKvirOOwmmcPpDujXBWno7rbE9BO8XRcPJXeyKSv6bBCaLN+cA
jfCK5F257Epzqauag+uqbrQVbkxuGAEHmuoVCPtKAM52nfnjU3k1nI2xXb8puzWQ
jyVv+JtTSSBWkHWntMRn7Tlln7FxIwnc43AvPyeYgJ66SyW9Mx7oA+Moh6pep9ic
9NICET/VuX2Dhgy3nxBaQL48yVu5Mn2yvcqZVkpv9eSXQUC/veRFhI5RxUN1ITCb
QNSti6GJA/LqZzzZ8iNfy+RDXveZFlJ+2Pa0ojAQ7WyxAfkcWMcGkVmgQQvRcSxK
29RWHXu1up1ioZglNHnjcDtnnUrgMviPWHHLJCRh/+KNGrQyy82obY3AiVzY/Ut0
3q7ZwgOilNF1ftJ55AwtiI651bGP0wvqFWrCeUdpkCkDa7bqfl4aJOmopJjMkPO4
kUGqtzfI6iID0olX8NB+xW8kUA2OY8OvvQrWRrwK+mm/HHWS5E30OOQP4+UO9cXz
5D8xh4a3LdrOV5zAQBNBcexFzg034VYGdOLcGyaZhUOQ7yovb3FlHTZHhnoFoBlf
g3YGI/GT1cErHilEYC86rxcgiYauVvEcY7zhHjGsWJ1xfXnZKOGySe7fSjBn3i5n
AWee/vkihU7SARMe4S60DDQTpFqgqp2sxqew537m4pdTHbbH4jA2aj1FLk1UxZro
02RpWGmVTZKIIp60z+G6/KMwvd6REihBwk8AkQeZgYheGR1MVTL1qgYtpxrGdAyu
Qr3LbzOvRVlYKF5vkwl9bAHbsFbbyRd6vkUUbqSslPP16++9zivHiGsAcu6RimzI
Z9xnuH1XA+CljIJ7wBp5n5DJipQV46UUf6yRFHlpYpSHOPIgo0zD1PLilEr0NlmZ
+X+sAWO029ejrdrluZHTq1VgyuCQYB/E1ZbN7VyUq7pceH+HPYdiuNqhhKluDfPS
78RLfRN1kTRLp/x2G+taRe1U1DokLmq7vJByzxechd1UhbjrHUXSN6ZrOzLLyKw6
8y+QscdCCtDrB35e4EIToF49wPrTIMcBCxCkefsqnOD6rcJwP3HfCs6A7zTop0VB
FmG7VYEjd19ThNmXx3X7bLtRFDQoyzx3eAEVJ4ubeBLKy+3m4auI+SI35qiNlExx
QRfUaE5nYPgpwHmuk5Vr3SHNW44oZbzonG08pBShdxJ/oriLTrAkiipkX6/Y6eST
qc0JAegqNFSoBlbzbTVtrAaZupcZO1EYdZc5AFBuBYRpntENa2W2t9ldgMOmRK1h
Xco6xev4p+8Bd0OeuUHE9e/8B5+DNHfpcWzjGcKeMUhrv/6WLSGq1My8HLDve0IY
QvzMbC+Bw9YksJt/QL+g9KTRT3qNOQ/sSJGb6MWKU64i/6a5EqRT449KHiPmX9nT
/Q3kEKyLlx5jdjZs62vedkSBDJkM3kddKzT7Fqzl6dw0mPr8ohThMU9qbdrRih0O
WUP8gMV7wkB7ijpU+GO2UBbAhV0WYHg7UFpwFygrvMIDSrcltP0PWpwUwrUdRObM
JP2F0BmUNZkSaO3D1JbPVhCrXyJI3QdOAqi2Hu/EQre4/pzmYyzpS0zCqA4UQ191
pwqbpr0UlSLAB9rLElco8qJ5VIVehLgXgzbHbzgKyFZk6ZWm33OHcB1pKWClx4pz
ChQlGOlYVKE5NaLev2WC3/hTogcvhRCLG8rV9Kg6HTCXy4jQLXbCJBPOHWahyruS
oBW9oFqvGn62d1eKRLbmpJl1/gWCfM4p+U1m921XNhkeveSPCGZoQV/VAUhkwnhG
f6glNzt5Da6NRvchQD0/Nf5kLUaL6wJXKwomRCHNhCG1kdL2e9ygmOb44hniaPjR
WWm7lyB2Uo3eaLUGSP5Dgo9Wp/e2y0+pxnG0/B4DXS3kBJOmkVGx888jXM+YKrbJ
UOVimdSamLQU2zyQBIQCnV0U0ROhcyROXj2eglP33j0VraUkUc98eYh4a4Y3IU+T
3LoKQsEtXXtdjgXcOI6y8UtG5k/hHWgw+e0YIv1M/VsadMVh345J5SWRAkeJKvG+
/t6a+id9hfE54RzQambLKiSG1a2BwhizrASq1s7SSZbPVh3u5rltD1A91/EV7+u/
3XmtvFu3BpPkP4RXdAXtagKuw+4gIXpMnW4GHNOVh+L0+RKJaP5w2PtTiz75E8M0
EXTOc3SJ93F/+AcRZqQTmz8Mwg72qBMue+xc2FxTsWojdokrgSak8W7s7s0FZGY7
n0Acl4Sewhia3h1DhXyde+jljc4MgsOLYzDmCJqqo1e8FpRDAgSSEOw2cqWMZHkC
SVjpxjr92M/FTI/7VcPivFYVoCl6800hrH10y3YbobZZyQdn/bY8YN0OLNcyDKVt
J3rmZDMErQhGEWDdBch2qlwNxZr5ymHADoVSk5lX2XsmStuh+iAtrCtLot0DYpgf
/oHhkRufmPcSk6KE5tJOD4JEBP/2hk7TzuZFTNwtjpUtYBQURgqr+NSpKx7OeO/c
2g+Gh/G5je2vA/8dUzDDMbF9vOdCHqEWcaagLua9G/zwYY/hqEaohvQ7VSNBFH0l
/K6ma9rUK67DsdcjbMpFowwuLRWsojDW70cFmwODNeJLoXrG7T9CWOoqL27KgBmQ
zogOM/RuADkxXJTeQDw2l4N0zxHxi6+rKjCrkF7SNHL71r6DnNK18gJ1rbzvxEK1
5pRb8Q+KctnFDcL20/xQQ811hqeOCe2p2YxlPT7aM3YIxY1doceaGF2WLDcCCusn
xWfpRvmgBLn7zYdBOYg8q7UnFiIjVBdaapto/bZmKwcKzC3W9o3U5O3oqFcYPCeD
eZxZx4cBgCb/NfD8XbzlvnaAEQ5/fAYwnNQwkjxozQ1aKiFap+1U98s3e47LDj4k
3a5UkjvSswJRqBqUWwg4s+b3qBu9mSmWRoOpNPf5UqqdcX2ov8qwMmiBqvBrbMUo
3VbceLLyeGTUBxDelMJBMofXOs+JIS/tURaJSAMLu3Pr74R8vitj6buesF6z+6L0
KmYHwxxsZ2dqX4Xr/jMi38FvV7nL2UnBp6pWTovIEJJdBZLoYlXDN9qypLYl0lPA
VryJX8tW11Sr4bkQVS4oqY8boMbEmVQ3mibj3xurH3O+JPuWl2RsFIaSAMO2iDF9
E7L1mmrBowKc6VVSmF62kMr65x/UDQrMdbwXkibv8QbuJCmQmdXAx6gWQhVyltNL
4x/uO7ST0DMVqs2X3miGs/vjUwcyQrdqJmsvT9WBReKAZBTVjqe0gCnxlafbkf3t
iiz4N6le4VUVCKxu3Y0JAOa+GPpoynxw0QKExkmGlMiSq6awFpKaP+UZEsIb9PK3
Hez1TNrTIYk8N7TS7iZL9eqgCWnAxZhOIOuin6FAV9Z8behzUfmbo3LI1U8kBBzp
x3tFi5KXftniZ2so296Gtk5+kPauEWVxUa5/XSbCnlxL/+roktgmWn3pWKL9iPQW
jT5wGTs9wmoj+4RXH+9VPxHMpB+NTwIMWuJ2bf5dTj3xfzPcallm4S0o6hl1NS6s
P8mJJDRHrlnM9dwKX+IJFeSRuLjm2dUa8s8fOy+yOsV8lN2fGhPAhQA5FDu3rC6x
wJ2a7cx37V/acHPm7fAw9Fx6hNiujycwZpbPOKQ6IAjrpj7bLqPPsCSpk8+Jhscv
CsL5UyiB7mrADbd7JSjJ7agebIQu/ge8bG3mySQ/BhHCgqEYni2HbTJv8t+y6wZM
/2fcaE8d7kYdDeyTN/dlU1vpLjCZn5IysJz6IskNK+xH0SX8DqVNgXEruvyCzVwR
XXSwdkHBSX3kJ0Z+P6Y/bACGvGURNMOwzCiHcsM1cdYQeQdI5HfenXAp44Jx82zz
4zW9iHD5MbKcnNgi/FKXGpGucOGfO4cgVkH/4a7+YAP0BmY1CYDjEHjm+xdaQUby
ASB5BOP/JYs5jcxYO5mZPWMNuqhxgnxJnEVYaeK/52Wkm4TDDRJ69hQobQypkn4t
8T5vq9FvE/C93HazzAM4sFF3JFdyOxGObl8yZ6JUB07trErLTlyimnvy0wy5XT4a
a2OHEZGp/1q8jFdniIIOJXOz9qHZm6QN6+OeTxTOJ7yOEs71kq8LbCj+ZhEWjeGd
KA5jU9P0Gn3ESsMhVX1gfqRUjtv/ZmdQVA3AzQUqL+QhqenWtf/7TMeSxtvUBxTm
UCYZ/VSlD8subGEFMTriciUmb7jcWlKvCoHj0/fNaz1OaLJYIvL2jFQr+bNQbu6u
gjMgUU6sLxu0GN0EGWAf0OZcZd5/aohxhtYBMFPrKaRKzaGKcq5epNrxtl5qbAL/
lEljvkElWWqIHulv+ZaGIYjvGu/wNhftptt4PhrpZ9PmaPaqJyCmZ2xEqsHW48ZG
cS1NCHN3+9hO3XJjor6UyBHvOMxCbc/edIvY8sIAckNrZNPPDIsjlBwunZj7DdLw
8tNzxocCuLIEIslk/lfibUXMwSKZVfmJyYQX5nQW7Tejm42LndZeaSjKdxG9QZFw
65uu/FtlznQLn2XgtBGy5xCDazdlAYB6NLNpSohuXvw4dEhjEIWi2VItiljwI1m6
E4fPPzr8PRnRyeLqfIAH2OezITOKof8bGDeWJto+m0IatBz0xQJ31VE4pikyl60S
pynX2OyGkMoFuG5YBlj1ySV+p2WO83MJx7FSP3hxSiL9EICuFIxxYT+56D5MqLx7
uDLSDzZfCT3uiLdjZ57QM+E2Otr6j49omrnaEHMDEo0V7lDT6qZngsL4mEuJkaks
uTIiTYGFaKQNCGpCaeiQjpHOOde0BorSpr2HqEjndxNLM3/yI6WDQi4NI3FDELgy
ewbABiCVj/E4SfKEMfsHddo/MPwrizmFHNmBoH5/aArx99BceR45cY6jwo2MZev0
yqFgfkGlmg2JFva13kCnsAbDMf6FPcAiHHHrGcYhjsHDjq8zs+m2eezZqCLSuOnq
7oHbBBUHHh6A8Zxc3eiRGkMkQcLV7emzRD1OV/N+GdjeTh/XFjKEDyHbpMcHZn//
UAGVFuK49vAAJBULRdkWVKqXPmTRkXgy4X1fbG/Gzo1+lDbGtAp/mJliRmJn02y6
Eo2WLwvI7SY7BL0hjQGOWi1MCNNU9OAtISkJke3w3vN3LWl4RH7sfhdcGK+qUtyC
EQCwexXWXVmkxRsLqfTRcYYcqnS36AhyJdNSF/knZ+fN5h9StlsjLzvDiZsR816y
YWOZGcsZ5+s1IiL8X6W7Jja9h//6fhHYPUzkpEEuip+7PgtAvP6tXkumSKEY5BMe
AagUQ6xUh/5VP+XvymYbm7+6/UzHrsJp6qZNfdhzSzEu2vWy4AfpchQq/IIzTQco
wXF8d2LarhO325Kql24l5Tn8ouoaqYU/L880SBV6it2J6wfx/HU9S4bVz1ARn7x7
7V25eIZn95RbAdLUcp299HjC2lJ3QSnw/PIiLjnRUKW4v1sq4zmBQBQK8C6xWq07
ovMThmdogT58SSNqPM95PN29YdNR/L++1vtmEbYvDvFYdBEVZxf1jXi7T9cg1Qiw
650gu8Apr1mikT8uOg8jJEjjqUoda9FY+yWARQoVn4y0nI19wqVDGgLe0WD3z3f9
K9SJxQfvEqa8RPiBrWkY+PcVv5IAZH7t3dVx9gSL26QF8q/1jQGfxLLYrRRBHpxa
AtiSmXWC/T2qz8cnIOB6wCx1kY/xdX3hQQZ3O7TejAzIJLCuaLIG+Y+Kgm7M/qx2
DGdxOcK4cAiqaYmKvx40AWH63WvrRKOA7gImFfT32GIrKj2/Z+5sMOAEEItVxhFb
tI2PMAbGeK04Be5sNw+wT5dXH5QYda/8HK1g/h8WN2B1fFaakHnEMMlruV/rTKtD
daZkffViJGCHLRNi/apfS08+w0KEHdLagyJUCFiMe28Y26+wtXiv6XXhQS3qMEBQ
HgR5+hXqrpQ2DwnGAVOMwYtxJPdIR8MvIG3Z3JHwpo9pULiLtftSK+tMrZcsWaKi
6sWzh+HhZX16jCQOLtnH9CzFofT/FvtgSj2BDmcBnWqCT76j/vDj0skWe4Azl2/2
G7DXeeW1Zxe2YP4Wyf2AY1L7OsUdeu0Ee1IVAKw/jV0QDXGyF6TpgBrC9lk41ATm
5l4r2tf2H3M9F2/N9LPL/IN5ENFkb99DudotmTNCzfT2sA4r0BKOuzbg5I/CffVC
0pW57fuke1tI3JH77lDx4j5j3+N7S7tjSkoi4d1+33QyJlHIRQcBBk9+NMAWgL/c
gny6wyZgkOcTJrsqjPzAmBLY7jbZnieCFPA353Lf0rNur0lWsyfXLBxOJnGnFWbh
mumr6F1XF6udIgdu1BMDdwXYcOxo/B4IgrVaSnQDKI6ZTo7fSpKnC/ncH261S1h1
cIdWOzsoqHnMJJ8clVO8KmyoNwMfNdU4dREeLEdTD4cW774mTVPXBxTdz6lvQvaV
KM+lowgJd87m3Ipicw5kQMBar1TJeWf2Un9J6FGxWf7yh4s5GaUg538038jgX0Pl
PM0ZEejrl+ObljeWCuuOMs2fudXIVBf4V8NgiaCNv0AVd1xcxHwsxUZqzB0pcgDf
03HtiFEJuK3Yo1JygkzaGfzTX0KSjf8PhUqsE9cuLiRDX2hzzWCuwDx/NjIN0Tar
4L8WCgwlwWtUiPzVNOdFA/070E9kEz0Wq21OJpb1i1IPSs/QC/EdHYbxh1DHarb4
Ja5VJeQn5ceo0Es2DYvvsM3C2A6Md4vK39YuqBdXg0yWVqqqIN3jTLADj49g30P7
9F/ib7/vDBVkZ/xowpCG1qDg11jg0QtDqbMHRtpm2oIqullt3W+jE6HyOEJCEByg
lM9MIveYUQLPVqRLm0DfrqTvQtA2oslgDSV+B/HxLjiCb3GKHabkIemNpmu+uNcT
tLqA7Ca7MwQkpiHtDCQakL1TVl8fAlDBMjEukalcu2FhHdiivju5Yp5cTS4aBQjZ
VQ+wRoNdbXe9GiMiiC/uzYvId2iUH2TN48FbP03jD9mklBH3HAkmPmz275mtPjbc
iFbhDmfrgwLch+HJTl8J8tl6lvfKRCVLNdOfPUGH2+H8aYDOAzfwIeFAT9slUK2J
JQADYb4iCmo6bZH2bNXx+WmZt3Fu41/vIBEY7Mjafm8yji7RBp10t5lyf1iYqkEI
TxGo403qNf/SKzoL/Ajghfe5bkQsQesSL1RbtL0WpKmb9Br2jweQyG7KJfvONW5l
gpZ56qM3aFot93zVpLc7UYZVNdxz2tUtAhTSrkQ/dOk8OzpnLVO8uASLfsWhMcSe
dVQRWCBIF0FY54MUE5nTl3ZKrab8BJm3n7RYDdQELXE4WC/Gwn7iztaHdyZ3ZLWh
B2n7TLUrGPs66VaPY8KtYqaILIjzSETQr+mgBoA3IgsGfzIUo7CHp5WYdQHXnsBz
wN8fc1jy/vEjyYwvwqBzn9RgYPdOYfNbEp9hemuvx3cG9cqzL1kWq/nAkGAvN9P2
b4uCsZ5zv2cXyoyOuDsZPmBqHW6hP6LHG5rSjg4Kr3WFxn7shQmccNS9kuMq9psF
S7HpMr8myjxY28C5elTJZ+y57vtJk23hGswhEgYaIXRRQMPRlOpqOQnzRJVj/2G4
QlftRRpnJXF28bpbFnoyvS3BlwJ0SQon4getj38nA2EM4BYaJaLiMvuritangmA1
KwOQIyd4Jj+/4hO/pIjylwjBlDupq1UF+nHPPZsjXRF+FkqURR7ga1tW3kZYGxDs
gCjUH1PveYiFSLWkPviB56tJuW5oZ5HBCo8sWTFuIEU0iy/96Eg2vaKlEf2Iw8GR
0Gfs3lebdydjR1hgyi9bO6SDo9iGqhWjgB0L5u2Xgl76iaMdSurQofn6AunkuDrS
dpsfdYpiW/SPBPEf84uWoJz8sAgbLb1rJxdeGjy7V+pY9+EArF4MYnRxzAv/BP07
102lJiAwBv/RK9Tw5OMs1wO0sLkXJrPRy43B6X0DJeTifMZyFyz7taJZEP+NFjxZ
U0Osgl0Sn1C1Lb+jRzsvVA1OoAuMT9zdr5gC5PY52UAs1+0kLfNhJkVFJ108WtbL
IE/6WPzD7M9sRt4ojZiFTccsZ7Wpvl07tVLAboZKHfjQMxv3Mrc3zOk9cwLOXsVH
9o0v4Ot4j/MBRWEVyeXI+62NUXUMDN/0sUf2Ma3JZ7k9TwpUJU/HRe43F9VBk+nq
Q/FJTb/wwM3Ddlxb4VDooNF75rh3iDQ9elKm5hNOTK/J6+/cxwfvLjc+hb1/3NZy
nzeCpWgyG9b+Kic9fA5lsgJ0/qnTmE96lgBKaTUrPbVo83jfzAG5rXUCJJ2Fpopb
/pEkS+TPRafiDSSxnND8ZnJ2e96kWNQbQvZP+Z4w6KMqpgGB/arRePHX3DQA/Hms
Zngf0CPj9KhBjXMdf/UAIHp3aytlbtJ73tLkAzkHAJ5iwuC2LjnEQR7mD6PsZXSp
92CJoHGwUkWF72E0TuoiFONMXbRb/ZqMEdy6cJhgCsYmY6gQSSzsjwUK5JrGa42I
iF7vFwoTYCR6kmp61rtV17a0yNQealA/AisglxM3bibe4XQsF9wJMVm7jFXwFV1h
NtMu+Cmu4hg+NBUoRKF8EJVRtO+bGHcR7ua5sC4btYSI/s+RWh/Jw5B7A5w9awSC
UmbOW9STXFHRSjSc/op2OWYushC4EtdTE8QmZBf8UvH3htH71iqVNnvCVsK55DCX
Wlsq6ppBnZOHsUCxfatK0wlYsnhkQlzEFt1XKdUF/naDrlld/h+nViQMtvbAFEUV
YFAz/9qx/IdgqIuLLapqKqgKw4ief2y/it1QKWaigIGfuHEhPJM1iK8bw/aG3u9D
TwALywBEXGJLw2jLvQB341E6E9mpWZld1cEXRzJHUJUFQSKigxgxiA9yv50ReWuF
Du0V+v6OqIrvm6NOiCh2lkMMeNBRYkJt3hJDxhZSvUs97EGUPnFt/J/kP7ewYhC/
yNZXPO+kqvcA/ov+8OoWivB4AylaU0KTr5JAk8dNdwlQ7d/FZj4h33pkwJH5WZNi
22Mhlea8RU8GC6RUfNqWt7QwF0Wl3YpnusqVsQqWFLqQXEQMFVz+IudJY+QFOD/J
YT5wFXgEc4/bbVsWCfNBgTvqr1po+kNZJm/CN+xyQvsANebJACuYQW6LuJqKLYY6
t66jaA0tc9UXiGjV3b6nh3RNMCSoZ5anpDVWdblEybJNwfV4tEje9fWun05AaEk5
vGF+Bd/8KW2meVsrVV3IibXHgkeledVNgSwpqZO5Sx1McjA1GPiXdcGZaSLUwnvD
x4Q/DsXUTrjQRN4vNCtqhk7V7rpZTbWJky0vZ64NLCuy8rugx8/LQ3xc15r40ufz
ERBm0E+p3sV6UVMA1tQt7kQmm+f6rPKV69t0hoxd8IOdlMyoPaGFcP8pB/KLft1o
etNYPDBFz7vG9YUSABpVscE7FHPCo/V/Pnxi0UO5VdWWR3krF0N5X9DK1wubCwZG
EHda0Up123Td0jxxbeOQaBsgXKew/w94ZLBtkx9usg8m3/McE0+m3PnPXcUv4TdO
grD8T3Wnx0V+6uG2o0qzFYGJgZSyNrfJwPiF8Jk9C8Vy4AavaXVkg7L+TGLHoOBg
Qs5HgD8LZFpAS0M5hlAtdED4E/wCExbMzMxDgLM6vq+1A97ifzaYjY1EWJ7O988y
09/gLu9jPDoisBfsf/tGuGrXomxn9MWh0+ycU1jZBS5RPNWtH+1K5O0qpw2xitdl
h2q39GbxFn4m7+CW1hkfQpPUgLGbvYS3CwT0awIOMQlPufceA3QEF0CgOjPt8lm2
a2UMBRXiTOZIhxvwy2iNemT6EPN0UQBXLDc09YvUaJw5EYas6yY27GgIl8/Lf2hb
9F0ZG9251WZrXpdJsjNZLyxuHRWHfS4Vqxx1XN2yuAJtd7LtywgjSGtidQ17mR15
rZSxdLN3Gs87HDZ0pqSsna0Lps1u41dO89CDeCcASRLpO5Y9JIPTSMYTfwMVi+Kc
T2YV9pKCbpmFJLo3JXK6wouyaWLHy8ehoZBjhkayjOVAsvehGe33qCM028sk0OX2
uRog1+LkmyWhQkMTO/ZQfFiq9YHHbLleuEddhsetTg2vT+9ioeYh+miy1SBPi/Ul
Bn3mTiL3Ftd+/I+Cj3IMGdmPxm91d8moxJE0VqamxhGl/XW9RVvMF2vxzstTGkn/
kM5NKWp3CTeTPbFUCtIuzhJYE1XdgUKtOLkpimEsiG85jtZIoGdWoE1PKH7hlk6A
Xh0rfsxE22AkJnUvlqo/vkaX5wFO44APmdi+HTb4ONBtkd2fNQ5mtCJkSXdtPHhh
vhno4F24WGsSpIPqSaP3K3at/Ou14toC4zUdnodGGqha1TwuSOMhFqw1pi5gTNBk
yPkeihEt4H6Ig55dQ+eNAPbl7nIKh2AoJ1jWMaaZjP+idlkfM5nWO/0eBbGgtvWT
t3vComWk3d8Nd0Id21OKhvnrKMRvYs6cliIRO9U+8cI4gn2Qj9zbE0VknGssI/gK
BPiPWl8+vofogAuIWoixfsqBICMw4f0LFZKAMOmVvQow3Dd0LgfqKYFb5ZtYjPTV
q8/P+SP4d1EKxIX2/xIFvPG018nWwCkRkp0E6TZJvrtOWVNvF2TYD9rhb0ZI5fcB
UYkCrNHPsueWvhRuIOS5oW7CJUjWk6EGIHJEgbUNFCGalUZdTQyg7yTduvct+BQK
D7G+BIYwqw25r3VxwhWHq60ucBQozTwR7xLRKTDVU7HlglQJtyG4+lw3F+cuG+3I
HrpVHMDjyIctLzFUvLP2MWVuI6jiwg6PeSjgEJRmwu96JTM94vm/KInLd+yCKYYD
6U1KL5lKNxGiS5SKkgW5LMviYRhxaJwad7HLPRp8GuC1OmFngl12A/Am26bKOLqe
el8eCp3Rmdc8zpRe6FXEDOOnZgO7Qfxvc7DqOdtqnkkRRi3TRiTEkiUl309xRNjk
H8AbjHE+EA99B1kq7QlPaMuMGtZjmBq783dGff3PGpX3Go1DHYpe0K4JDaIyloZA
v/ZtclaQRl9u+EhWsJU4HoBspyYJPHr9mqrtfW2VVR2uxMs6+Vhf32M3mSTq6XAK
NYtzUpote+9EgOmJ5R6woa8/Ti8DiC/miTyC25OLQDiGSvc2/n4GcwGLBBnVt2QJ
5HINsGFK8dv8cUXhlFCj/7THfwBCz7NvwYR4tm05LyFgNWT9lbH72N8OrUz5qxpc
id3RcqrWhpkcjWH9HnEOt/vqkB4888EOxCm8aAWkCKHWAA19kKpr6W9+hs7x28vK
Wtuhwrlze+ioCcKa2GT6uv6UvjrCehnf233vnAXc35+mrsjmCTvQ3v6gaRMucSzK
EHvbkYG5uMf4lUogPayXkUcZ+0dPDDBwaq0dDA2rh8amNn/o8rXKVe5JJtCJLmBr
ld8itfUp7WcIgilQHFQV9IMLtzQtTR2KNNPXqZH29ivezTCpqby1iS28rLju7dx0
aHheB+3LtSQoeymL/VUBgpAjAa5hncuzx+vwVOie7dOOqC8rVTmfSb7ClkCtuUmY
uzNxjgH/ngfFyTxVhcI9h7KDmbYeQYu8jmhzoJ8PddThQrzxptu7/xFERCRIXIfB
GeUbpkwOVhSVNCqv59+D5HKD6Ko+cVl0EdRIZPAkQIoDTs5JXbroL057OGxfkn+3
zY1C5E6R5wD5/sYFnA97MKRfYZvMMsI8mo2c4arbDm53Xjj56hUmwqf0rS6Js8+5
csazOhdevAdNfKkPCkIqMbiuwVHZhRC8lSaKCdWoar9G8LmTKCGQ66h57Srl4Yra
CNJXd7teqvAdkMEpZTxfkn215MOakhSpILVTl9cnkWL9eNrer/l3jW+hD8pv0D/M
MvNYMwP1sU+qeAY9lRh/CL7elrV2Eq8xqm3DNiG0id09AanOuB/4sXaWddJ6f72e
9sNGiYnMNu8jvBSsexu63iNhfBtlNb17CTPPgpt4lsvKfATw13pLkqNP0GNwt105
8lHW+Cyq+VIM1FolftHim943FLKN6y640N1uNJ3/Hx4/feitBpdz/b+LdTY0mDg/
zonLrDeFUlQrg0mmhywNeZYsOB/ubmLsiFML9ydXh+ypN57PR3d8MxDE/IUUAnnt
ek6S0wjcWPlsuiOAfFoOOqIiPddxE/KTOg4Y8wbs7cOYjAZ/zoLO+XJCnV1XHtIn
wPMYjDHSg70MGdqNNmrpFLYGvVBAcWKLpgkXQjAoqORbV6J5JVi90/iNMPn36zk8
Ub5oo7tCqHRKa7FxBitZRNIe9Ve9bziQtAEm3bKc2R0J7J2LaVOc27LFTeNu+rNb
tjgI0YLPzkm0/n0q7U1bBnaZgbUgZcAqzh++RoCQ+qpyWsu/AedrL5et378rKJpu
3r6c9i7uRCxuSTlShvxtq2EupsQH1Pb5NdTpOlOSyK3VhZ3n7Wq55nPXjsTGVT0X
9IgIvj2RN5AvEG9P7sJEHRccofGYbvukf+cIsFjydDzNOMq8np+we6Gv2AfipJHt
12hxU7y3OiKvgjDjk93mJozWeJVaxSvFw+31tC5XVudLtmKf6XClqSDYYPWH2p5y
uoyDruPPDHPuUH8wIZTlBIWhTFgvolchoyWjrPLBWbLvJJgcOk0PsKHmoEtm7hdD
YIBAV+398LmjCoC1ywaqCtfyL2A3hOqH598I3I6/SC/frXy1W+C/s1ZjkREyXeux
qkGBkqO63Qp0euGR6+oiXaCUuzRvcr+l3JAKZmABMVFYdkbGtdLB1gqSq9/a5KTR
Xxtmg8USK19J+5pG+tWNnXOP10URED3SCP7eYSdDH68Ze36iPkq9Wc4tDpBEbU1A
KS6sF4X5eoHuhIbHT35vJJjDSAUf8bhKrVnqoqalFxI1c2dZHemecZ/fu7KKb0Tx
SMqkSDx5hgYoRJhKCxMWvUSme8eyjc30iDkaBrKCww92VCyhlXWFhstCuZ0/pEsC
2PmeTufe4miKMHK0puJ5tA9pefc+fNXdedidEnRmeF5JMin0uuXdkTjwMJpo3Vpx
FmvThTCJNGUkPiEFZT35dG1YKHnXZrG/r5kt8L7aeho3BGWzLE8uvErlwryJQqm5
5MCUv6FsgyqcW44N5lrutKRxrCT5twGzHf4sXOHKeVPdYX8GATF/V+ZxfcDD9ffO
PdlB9x8BOmNFkpcRKRLr8iVTaV2Bj6fWx4ftr3QAshGnyI4/jmiOK75S9QOQMnj4
IgHQwFB4bl1ugV/BilwitF3Vo5aTApIFAIBQxNZubfCgEx+JnERCqMKDo7AW+v+4
lB447HP2UW4zTGpZCsFkZ0rpnJ0w3LYFR/JQwChQER31Dd+a/i2fxB7V7W44e9U6
MX7ZH1SFFGp4SQBRCCzM5uH4kpntK21ZwzlKuAw8VQTbSWp5v9UXlwovtRM2bCpB
4Bfq62nlAhZnoB5ODgP804n3Kb0h7Ddq7Q2mg6gLXwgb4a7snT4A3RNLOgu/QhUN
zNsTRYR8G1jH+TN79751dVkufFWDXE717yeb6RVeN45J50HMtzfv5zc08JvzgrMb
LGZrRUVVNw+0BbQQcjGoBjoIksUjiPSBJ/r/7SiljzweCgMW3fWpGG5UHcWJJfgD
qdqN9sEl/+boB163+uW+mu4Iy8Es79qKARH8ZZoAdeUAlKrNKxUJZdN44LWxbTN2
TDPsR2hC9g6DP5LM7MPya7UX90WhmTsbdAMHfAFwkFs6JB2bnNSgG34mGYDiVN93
TY2wxZ1vkjx2nJsZFyu4jMDAS+MukeMv1d9xvtZaAI9+C5PSgBhl4khtWzLN+VA1
G1wjCODkiKBpQtaYyLEMrMmQY93M7nhow6bg+awtBC/Na4tUH7cS8SybKeUItpAf
hkMhX9ji+xEq5Lhl+6nOmWVsSJ8AAfasFmiE2nJTHMxMOz6lZkP9/fKkzMbbqxKl
gtdU+MAMjxjz/bUNuRvoe2rYinxD0edNAZTJjBLd/mVQuXtaqcBMPRT/P6iOXEXJ
OfHIhVANUu2gtzZF4EJG3LPSOWeqLNqaad3o7n9X8kPM/t4WFUlWQUFhLeR4m4kq
nLG0aaVDxcdnA1/2+rxEKsym+Xsw6PRdOBLU5wYZqzV6pAHe6VO0HHL9MPT2R5id
zUqpKzU/XQwFqiiM4i6QK7H1cACi8tn5W3z1qTGQ1kcNRaoHMrT78dOAm5bzVGpL
cD2Dp1X2CdfaDcTaMlBTQt9Por0Eigb/tcYLdnhuVt+PRqzRRJUFm2pdaXNL76iE
LST19JQ0ZvULGjFLeIGL1x2mlj4cMC+1ARz2U0xdO9GmiMqbXVOFldGKBMeugO25
SFj6CZCHA4pB1vnU/DPdjIWZ60yNz3qJZvsaUWuWj7xPMmtWKlf7I9veBl4OMjcE
ee2vE73cZvj+qKp/Ec4wbLoKdQ6rJPuL8uKC5sOvXa2Az1pSvAtmASG1QYGawHSX
3Wr4SmTO6J0zH0073kbigKG5JcxK7hTanVJ5WFgUYO7rKXXFZSPBiPSbj/DhSpqy
VAxWPqaXTOerC8iYmoeGEj0ql83HcJBWe2Ml9/87bMn7aPBVSD5iz7uYR+wR+WUi
3gOez45oDgzPTQQ/xlFndz/098tZp3o9wc5bY6EddIg8vA05q7EHuSFA3wFOMAWO
bVRHiBkmez+DYvafaYbNr+DcIR5SjA3qOM11tap58aaZfKPQRjVEUCarB9rwpAiB
YjB/J2fgCMr45MjHkfso0Z+J+CNcBI1dFyYQhUVLHATBHDBYTZac122qz8WFcjZH
p44jrBnIAxjTRbjpJmEUWFUtpzVl9o7W9wsWaI6BtGQF+YymG/6WjmETJRFLw/rT
rBalTJ4m4/TZyde7RJ/ovmAs19M1+YaC9GOxtKjYkXan51e6kFpfH7gsB8uQ6IbN
uy81OG1KFwvhM0rEwXROnLRzZJi4IAbTKmkVO/KRLLDxksXKmMj9uBcq9JaP/ktE
sfW/CnVA+bf3VMxQHJpoKyefLxhWnJaTKpv7FUON1fXe/6dalkFuXZ9CWKe6m9Uj
ycm8xkUWyfHpnaJvvSwBclj+wOke/BvzrPo/x8UH8C9hBrtwzLAjEg5OP8rMhQMC
3tVDLJXxO7tzlGmNADvAKKhkCYIUanLc7uE9IaGUpwVvo+/lAuUx+7VG9p5vbxDp
uDw+8iNpRaiSXmsMUoC0F2BAddbVo+9PGvRSvsUgcvfkUcjDgVgRhT+brx1jj29g
d/MUrfGS6dklfNV/0aL4Lp3ts4ZCXdGh/J3NJBYiJZrL3Bn/EwWCYxXwuvh6UDRw
3PbUcnchNWJuQkT4ap9/W3eiJMkxEzRe0KkEq+vG8AZoyIA65QEY/9R3ECD6hU6q
gXMGO6jo5M2Iro8GEGNlCgKCREBan+Na8ctfn9bwDxiEv+mkXR9FfFJYL66DL+AC
6PZUTV5fMTXY68aHpeTO9JdPi4+88bQVR1nSJzB5qb9EjgnceqtSqk2DcRzv1qAj
Qm9RFEvhWm3GghXe518PU9icg7u0ocWuTRRXbqAeYvCxEfJFrua888pndYbuUIv/
+YvFZB6hFwSGAoY038qnantwGhGncOl0pEOdAC/4pKucisLqq3NCrNFvT19JtSiP
8+9LaUgkpG65K72MhNqUw4MxVPc2y5EJjDCR6qUpfKz+0BKzxt4UQaahwVjn6D2N
fngW8Zee4OWvAWUpdL7SnBUyd/FVlroKKprNDayFqKsVCrHk1KRxgkk0FFd0aF5m
AWAigmV4jKVo0Wjo1hqcrLJWOsZFqSCQ0eHi+fWrr13CZTzJZz+Q9Chv0xIHB4z9
Wta1FqTj0u/rTUA2VLku5SH6Ex/XxNy92sCNr1dyuZ4/aUpro/sH/MBGAjfOF+Cw
JCKy8NAmm888zlCUvp+KNwe79d5vO78uD7ixD8UYjoxEguSJTjbYzK7AF57Yrtnc
wpUioOI8NkhW6O5rjo5BnhsOeVcsfvMPLRXBRKdWyLyjx6kFV/dspRgNfcqPzyLJ
vpR61goh5+MgckX5ykiCtndgng46a6l0rLfYjOde6X45sRNyfUNVf6tbwK/iI2jb
WtlSkIEJJG1fxWO2HbQb0A5qJEzasdeaeQVtozJ4mrN8Dy4w94RMs3UZ+IiasSsR
ybInYcLELfnHo7bPCq00SQwcRuy0K4ky3J69c7pC5yOeUaOI1MNhpnsbod38dOYf
1pPn78tfzjFWTCIR6gHaEzOC/YLawExHiN9Hu0ddgubWg7WkgKWnK3lBFvEvpvFu
IUYJvfFbTyDzvo08qxPuqW6ED7vrPszZSf+Pt/zuUW8lhvBxqLXII6g+R6MphS06
s2SiTkFwKpssZx9tP/jria72bfzDSHzmkv9tKHrwXrQZNetS57r5E0IEGpVCfb/C
/N0/qMGUO+zxXzhPxpOv3pvjpwhtTzZ/r58UzwCP+JcsqwlSRNRz6JrX+f5QKdkG
UZxKd2VFyJy+12QA89qIuGpZk/QyDJRILVQDkvTttUWzKU7wA8denVweih27EPnV
ERdsQj6+t/977yTuYQeINrbU19nbg0Uw7JhOjNO8fFv2DHH5iwmzKU4MTSRwp4Jt
yUgWOTSwzhaqIT9dvqP/gQexOhycFDiSX3wym+A0GopZvY/dgy/OevJfAZJzGKeR
U9wHnyETjC0nocgu75hA4Nd8LjoH0f9IRZfftT3kXnb0IzAayNrAXhvRfti3MyUB
BeR3S09E0MIEELyWsyAVI3FlA9dbKN3MXdsXvWd2nyli4pH1VZuGFiAiaezvwOZV
tuutRx/E256bQGuKXhU+KywKjmiLKjnsbpTFRKGW+g67w/er1iwA9MPVjAINGocu
ody2ZLreGi+y6G5OWCrC9yVW7rpYslVRaYEthi2f3PQ4RU/0rbaI7a1lIxaxmbTA
xnSiU9+hyz0HBKUy2OaXemrKYPCyOJraqu2KNFx0x8ALmYcGx1TLWMNPY/2s6xAh
BCAjMnCMi7Q8I1IE5oO7j9knyKceaZybJrw20fq/Su8G2pkMDkpJ/HklR4S4Xc2s
zSjTor7pcmInUL3KzfZpMTJOEGIoZyRjignHyOk9f2DCa10aUHEdl1BkXnqNWtha
r6TNeo4Ij6NB7VVNKdEBi+4hkIZCx6Zjl96j1wNzwq8xBCgmm3E/p1q2qhNtrVWw
f/26xofwLKc5zj9yWBGDu+xwZ9ej4LnxpBj14IACwHSF5nmbZH92yR3CuDhEUvNk
gI8hZq+NpzuFnK39w4g2nW0U+yQUIgqueIhXI9yfHFfhH0gW2RlJ6pTqNklSEtk5
oIsl67oLaSpnFJ8aEV+eL6k5vhbUor76lLW8Z7pUvIgVMl47yaH/tlAhcTdioTb7
XwQByIh6tsLKM4TcrjSouD2iZN5SEa2O8sNTJF0C/FbzFlYIzFE8LkKdcnxVwWBk
qMk9VwUcHEf6FkTdADEP8Sa/Y47QOATbJUvJK0oDsI5bqD5N1vMtoulDy4aAFnsi
TeGt+h7/zDaOqcYn3ATAJYi10MSZ0iAHlvaxc25WYKWTDrBGxmO0A8/85FnKJDqF
Twc7xnnPtHKwuAYs10RL0M0Ga0DPqdyCJgArRNL27egPTUH7wqcSmyEAKM9A41tp
OiQw5WTz0wczvkoN3CqxPSRbjyyG6vdRwhf2lZTxkum73mErDZeTXT57mRsjy/gy
L1kUHbUsaRMxLJjMoKa2J8IUshvNAVK7b9U3FHzSOlJPLtNpis4HZT3qR7CoVN+N
DH1W0fVXCi+PTo70sMPW5HAuv2pUy9MPDAIFvMg8luN3CovIlG+Y06tdXWB6E/96
Mb8ZICZI7dbPfGuN0xmI+Dc67dLeaLQC3ap9BCXABPdmCdENSdL/3YIQobRqOGNb
gXzYh9YsMnzWsldCI3mtFIegaSimm4wCWLo3N4q7z8DVhF5ptTAjbDqT3DR0IDTw
SuVNeoRJu9ilIRayCjDgMwmtLQT7hgvbalV/zqgYPtGFTAKqJlKUW7Of24h66jih
b1JL9y6Jmk05PKOcP/YgIVqqwMQ0B4G4Ri6oXhW/c3PPvKNzmIkoCF6EmEAzBM99
M+m0HYKJudbIE9ujLhHHiFf/xv2eIZwIIC1Joi+IKKFVrPdx89hZR047UNs3rTyS
T9F3O7qhukKIJ3X9hMy5ffDBOMBRhCg9FQrwXEJS8XtbbT4RgtyVPumVdxE4R6TG
yNsjS3XAYBkTN/6qOwiR9Z3SbGXk3wDvq5obZw4gwcR/D8whdO4dhmADxvXeqHFF
bYM37chMBu87AoqxiqDK7Tzqwi9cNHYM6WKREanOqpTwKkTExN/FMycEtPCApHj7
OGKNvAozqxJU15+2PCDQ2X11vLGd0D3LrxYrCjTEoHJkH9QQ2wIyZw8SUdLGCS9X
+IF7rz/ZnXZghsaInhCKpWDD8MYyBPBSygqOgn4j/YkK1PkQyIlzKX5awBsPEfGw
FGnY9+1+eiY6douN6lBpHkAYp9l6PKbx1IoTaqWTmL90xdja9rVJnizPenK6uj4P
m9khDvvmOmolEoLp+IaWkQ2fYbgOs1eIN0XFij3nm6FvlCPQCU3E1L7ECudKY4D8
AeDIxNIsXMP/IFexnuLNIviGQWWfCFXkRQh67gwi2aNaacqR5q0Ei1Lx+qqXM/iU
Q8a61kh0aRw9buAPNF7zifhGey5+ywnxPI3XLDDEGM4Y6T8PVtaw2Y+cN4z1vVUE
UoqCWUl2WiGoEl5wNu4MtaVP3JZ9kOVdDaAfIj4OCekgo38GS84Zp+YwmKZA029b
1JGmLhp8+TewmRqgnTyoOEVKlNtWgn+7vg/ijIuFWtF5KAP/lj3Lq3yfEtYcmvmI
X2Gs51J+A0H4+eVJChy/G5e3NyVqXIifGh/UFdTnPirxSlA3Hh6GM34dWsIGJQ/+
BIxhfsee10Jix4cwCsgUK27lznRIeHUqcSqWeWbIas70yv1pr3LOIZ8lD9MRUQKF
oy5wz6HBmjmB/8H9e64nRU6PsldgWSTqmOLVMo9FrZafkUP+lU0+l0T/eBxIgGbB
2t58WbCFiewseLru8o4FOZa+5CHoiBZmYD1OmDQsnlrs9wQTeSS7cG1eW99jHOZy
IL+ZNsfSjcmNc1ByxiwKCmdwZTgERkHE1DW4LigqxwcOpCMudW1RxvyFHoFFx80a
Ybb1tGOg6sYW9er4tBDT0DNlvTLUCK2Rcu2toaTOURsKvaJ4+JEh8kT8wGXQBf1i
4Hr7SLmw4lT2RlN+HYCvYw1D0OuBj+I+WN1Hn8YmCgERhWZOQcJSQ/jzz3CM5fGL
LZ+HE9tNAz/pcZfCBIGxG2jLKDC9dFeINHjj4zdwKZ+hNWjsytiKjo+HPjNaA4MX
TW/1OMD4QkoBXVJ7HvW6HdG/L/425JhxfC1Tie9My0Sy06QmFnhlke7pEBOKsI7R
EiLExxm9lBzKGExJgZSbNx4vlwbBcPheOx1ubaqrEJFcs3ns0cXhMvi7XILoIw2+
/M5FUZUo/lOePbuxcgRciGRyxWmyDuR8AVyjWeuE1BkbwrtqKee89vD1R+KtqXFE
oF9kVQtVw4pYYOqXZk92rlXNiBe1nbjJy0b3EEczzjiE4vYWeJDS+ED9vbLmkVfY
spgm5gt2tsOhJDc47sn4VrfgirycVmkWz6IN/fRJdgz9/RjlCbZk9ZdNEht5D9ov
3JSfm1B1cwNGMZRP4pxwgArhn/AKR67EZj6c2iRYDBY0nptghZ5Hzee5MpQgOqMK
sRzo1EjLQmamiFgAX3uHqnCyhw31gORPuPLcvvvrE19jdNyYxJigNjgkJ5RBRLER
qE/tP0qqcFucdJYuhK6J7i13zIqEJnhWUhU0WVjbOupOmgICl1J2Go6d34JSQ/Df
TPBj32041T3oNA2g6Qo4qAevwLsGQiiuR81fvylCDOHjiVu4PIL+vnZ5qBLIy/Ad
kP/y69mz9F/0lhhoscjWhxD6xcDIubRmiHur9xCQ35InQM0vrT29do6o45ho92NQ
XqP3+tKNPRIQ7z2rkyQfcowjhx9UhEjpitWg81+USCD3SOrG7vYrjM6m71CU5bOR
7vEIwaHplVwAOzp769g82Ls6vGA3nb4navkjSKpUowAmPOLPovufLmQfWRSbnNMX
hup9e5uUENyLCNN4J6Ro59AstlTIRfaxnNKgb/UrjH58yxte5Uy9+nqStCaSOHsp
kTM0fnOMDdAcrp6FIpTJf2mUQGH5UePgBMEL/DY73qmY2ANvZQPKWl4doBZRua1n
Gs/+NHNxE2zuALfMUMVcNf/I11tmJJjf/vupJSaeiU3mrFliyw0tgO6X8QRazPgW
Hl8rS8LoSxpfvfTWzdWU+Vn+83AKn4BM9MSoepkqWdeqGWsZOrZbvMuJO5QNyGmd
PlRQ2SuDoEdO8b3J/2oWYp7LnrLGsoRVcmFfhIaBd1iG0fz3BO5Vdls9TtFvUUmh
CmCgPzip1LAgkd7664/wCSKqo87Iw7+gb1otFw3Q1QfK0e1F/VieQfE2KtbnFS3J
x9/LpxKYSWf0GHo7iHN71huIGlE0bH1MSUu7DBMjGvcqKKJc4/q6q3+U9cRo2+7w
PAtTI5cvq/ctvIMbR6c/aTDjLLVr9CP7jUAjE1Icd483jXzUiB3KPlLvAwdDiBpL
zWSqA6RYBPvMloFnVf95HPxr0bbe2TpE+QdcgZ4+zhadKJtWBlkkXrcIuGhwb3/i
w+LjcEe/sWLONIJtprWUx51LIWZ+RhVYCUa4LzYq9kGHkLdUE85vJGtJCWWsHpGH
3c/L086GV2rHaPZQ1tOf6XrFv8cwvrcrjaLcwy18Vx3qWRroj2SeRz7yH+qTMN72
Zm2ovwbHFSrIRIWOh3ikUEmPnEUK71n6hB1pqROZScOniaGhLI2zndL2nxLum7Sk
RnJCnMpuuiiZmQz8IIgj0QCyA21+1rGuy5PkMg6SfspYvSnsn18IfCdYWuzUTHhj
RDwrz1VPq8fMOAuGgfh/IxBJKZHzrhOrBMIxQiscQ/Cs1+RDKFV79M73x4VqcGvf
Oei8kugMtmcFP7JzTJLAvq/Q7cBdSCnBevN7DMWiBWcXhKldwyp38OmTBZFwzYKz
Slrx301Tb40Xv4qnDl/YMhXQ7lFb6zROajKI3DkFKGJSLy0265FEJ12/xT5rI0NM
d51zMheo/hf2Gz32C4Xy8UH/pn4gogCaz4fbFlF1IimEBjgiMQR/uF/3R8aNOx95
x4s9UVNWEIdI/3uPtoV4EynRjAVunY1K5fTpgEnQ2Ib0sp1gp+lm81RIfUNZCKFt
crNaiq3CCv7IB61YdRgioa7Jm9U5um+TbPHS/bBNBRJLEOY3eY94OA0o4NP+L6jd
pICdqdqUXuzXNFCNLpIoQAcsseb1xTtzS6fMsIKR0jDcZsrvjNl63YHSWkO6KlPz
2wazqXEgN1BYceVuOnVMawdGvMGKRNFIhtcq0VRHLjrtDmR/KT3CaZXAk8blwzcy
+eVmRrrSVou7PJU9JZqqnrX8SQYOKh7ZTrrc+eCTxHuavGBu6XyjdGx5UkaaLEBD
0MnuwjgveYVmBo0g0MnxbgJ8wSa+I1vgjvQ3nwQ376mqwyL0U20FPSCIPQUrNyv2
Bq5B1xWllE4d6w+DiIJmMxGLWpTaJdWxsABlCFN76ioxMxIVYu0lOqckvLqKjeXb
Gebw+QnvVKtZPfF+3i+GiB2RFB0mwAQt6h3s3ZVWqxQ43gilCKJ6lT6DUmoRUsr/
NRjodcZhE9Hpkq7wZYch7HV55mL8WYvU/b5SuRMhAqVaFUKyabF+y4Yb0WAeI2r6
2SMHTIg2h/6YDUWTaNq1PDkzrZIBJsOjDMIB5lzzkrkmEY/EfsQvSd/og4NZZeoE
zVdhng5SzM+k6zL1en4e0c9P4gMv1SrEEht8hHB656kPBBfNbYB0bLtPjn76a583
vPy6GD6JI0cBKUUFycDaVKIs2g96paQyROc6U1ArVwxQSBL49m/f8xDzCeYNen9V
j+1fcfvHUzZXLJz+8Lp38dVPhHdlhQs2+WFetHs+8kDjBk0gI3w7sW8v6YIEduPE
x/6GFuH9FYHO+zV0g86ChE2814U7KY+Vff6+Dg2/QEa81hgfJC9U2K3vlDGIEvUp
ax6pj9utCSxQop9NmQxF0TkG8mUxolIMIKTOwU//84mQA3d4Hg8XvSpWuZ9ldqPi
NKGgdV6yWuNRHQ/QP1tjRyakuafXNPuZqMjX4faTS6E0q8I7FuIHuieod/2tLNug
xVcGErOcu4ubtrvxZyQe027aWvQV1NUhrO2695jgTH80WHSCYpyyMK/Ido48Rv2A
oS9Y8pbkg/2oiqJwn1OpGxqIFxOZm4UeDkJ51/rVfdqiMvP2W0eH1qBbcGXg9WSF
MbuuVwiEmmFSaY1biSAQIJaaz8CTnZQbjS8iOQDbKlFd8FFVMV/i2xPUJpC+iUgI
XabLAd3Q/kb2IYSmbWQoa1GCm/RmoTxCOxTmicER47Zz+VVEraJS0VkLZCthOwA0
5yz6iVBz0VzUjqOHx4MdUJMtylFVsaGrVgpdF4KH6T490xFeiBlxKJ4xlrrEDsWb
Rlh39OEh3Z8lCA7p7/YgFdM2vCjC032sSd0pOgn1OxB3otFLrE28qKtRJ5/HZKoz
uDURHSHr0mQ44jJQXdCCsVz0stnn/YfmJriy4EJFhl4ApBKh1BPHrS+zHtEX+zIf
8lsdwgNLTygY1JjJhfuRIKhyoKYwN5totmnPJHn1Z26So5sVGoifux3Qb75xM1J+
Wja+V4q6VnE3sn5Ep93rKoOjIf/hNXQVA+HkkjslRxhp62Y80FASAi9b+Cxd5p+6
lthUvKefM3+nq/u6DOfIgdcHmILiZLSVZ9FxNoHRmGk+l8zukpnLcXB6MgqUzrib
Xj+acTuBv2AgeNJB2LC9qTZUlsq5hJaGEwjZJ3AOhERFiHdKZ1mPFf82q+kKhGvR
FWCUDnjW/3ihWZ3/7akmMH4EZm1uuXEnoZ++DwaPNVUlXXx8SgwibFZt/NcgDNs1
PQhAfuF4ZBpvzXGoi4MNUYo504Y9368yn/b4OTk2vZbTZI4dBRnXJ6/kvgbJ60Si
Ys5G8nOdMrLcSpVfQB6+kDrNXovQ0R5QHsVtCR60bantaPDgy8V3ffCrEj0yD3f3
DyPGqpwZxDl7Ft1JAfd+/AHyrTzPUiIGB6YPAsvk3JFpBIo/8nxvvMlmTcxmhACf
4Rg7yVOgkk0kUfagrCbuAS4EsAExbOjYavWCM9bey/z6lqC6acHVyY4izcwyB/tu
ijA4+sI5sqAaCNFztwApeco9GL2LGQXMPbXyQ192Xsj7oXkbWpreYl0YlWQVcoxR
y/Izu4OFZJYBDmrm7SnMcLQ8oxLfkMMbEd9CyT+HZwm9Yuelt5XxT5JEvCYwej5X
tr18dbArLPHocbEgT2ghgWav9MtegY8wzahMxpj6z2VTELtD9R4QmWghjNZ7Wqh+
23TcmyNr5fonIOTUD9DrL1gDoaCeQZZIaaHvh0x+I2o2cAcJqAb1tq+Qmb16BZiF
UxeNb/PYXAEFO1E7kP8dP9c7wPRuXvR536zDBQouuE48VdX9aUWWe+hlWE6D7BDk
C1/ilVwCr8Rt5yN9Q4Pl0vE0pnZ5RTO2bvWwEzTBcUm+j4+mEGvSmOl7nMTljdGw
d1cBtES5IXrE65fvOOnqpRMe/eNR4jZKrIWWGs+dcwlu3nqIaSBOh97HLC+nFmQj
81rcWLZRYN9Qzy2XqUEea5Ylnj4iSYu0i7ZU3ghXbKLb12KS3GxACvYuTkuEBxa5
DSnoPQOFTtZShERzoj2nZfEjq1ztBnNWVAptTgxPQnSwIJoahqll0bpDizAMpzpm
owS5l01Xib+UjJYzEGeyfJ1EELnu1p+mFk6a5RPglymQrFSmdLQLGKE/1SU5S/bl
4kYhgoxB4RCbqfWab7Ri2iSut//GWI2iStZXZIHY1UEOaY3dAplGJxccMTewgLxg
QBXOKEOc5FcDZzxwEEQbpbojykFYjuLuyenqYMoXQ19Y1P7xbYFaHV5KPYxnk7MY
a3jHAR7XcZno3HdcY8goWJT3nbNzOJIViFrJwrA1j/411S2zWZXZUg8YwbTX7tsM
2cbw7j/W2+1pyGCDi/0hwfsAwu7DjCXLs2qNT4duiL+wBm6kgRzo5nv3NiYOXIKN
hLDy9CoO9nPjP/Mz+5etEK5WrW8t+26oxBpFBwdOQSlvZYPAQjdBni32cYJFGSip
CkdHkum81orMkpZU/yAisVXoEFERM2i8DGCvGKItsXXHzxubjaWr+3zGBbT2rRn3
5UCZyOxaG4lUHOVYu4ansxG+U2xG/gyxec3kx8pYeIjMTcl6ZmZBK98iPojhDL0E
JHR0WNa9nvPpyRWcrc7vVh6UF+4k5qiNOdkAZb+OLodhOjN5YbLHZFBhSoRtCdNQ
Gu3Y+FOZDikVX49DqwcwLDEAQKue10kgZzH9tgDXdZLyQNIrYKCuJkMntZm6VdtG
c/4CAU5qpZfOK8Nv2Z2VK4QP1bpYwAfZ5wC9BypvcVL3TjXY2PC4EAS26vIHv5th
qtsNH7Qx6XI4fsXBmUtq0RDrVVmECEDXQx9m6NZxpQJe6OFuqOwhelshq34PldMa
nIzFs8tRgfcKZs5/unDsZfNNxj2LIOfLN7TfMx+eYUsIGf+z8ijG+gLbvZcgiOt7
j3ndfLDqUmc670zZgO+OoIpE0v0e/BZUq/kDsKJP6Isjot7gDoOoAcvHhHQeLpR+
uqjfn5kVkv7mxXCm/BiXWjzClu8FafxMIkFyMhlem4L4yXx7bmOqjDFEUlLo4OIH
e+Wf3Nv1fiJeA6+cpKp/LOBfqaYFUjx5lGv+EJdLdGvsB0hlCORraJAXrgb2kYOk
x1Bp5MMsM1a59Wj0J3Wul9WvS2KydE/byac2CzeXXkODgh3PUH63hFyyU4Z0277d
FkguAVKk77fBIn0LTM1bT10Bl/GyAGyCGcTiX6Ni8m9Ey0+NDGZOQ7afJO/+hFIh
MCYYv8MH2+nMhRWqEQB3NmLxjWQTfmupidQDq/Ly9qWjFDyzIwruxs+sMbYwCG2Y
3QeGzRjrhAgbTEYoCji3btDuq5MgRK0nRbLc4GiPfm72gMvYLAjPHNp2pnp+VMbZ
660DgRZYItfQXHurQieHB+SFFPMTOGBGLb12DydZnOjxll0ChVs9SUaDZTSges3C
rDT4unEU1MmqOL6+lfyTZKmNqmrhs3UHj/qz08TSutmTmh7KCTl5uaMcMdFxWuVu
nofy4KqllG2hBkNceKi1dKqr4qCPi1+75CKguxBz2RccObTBlUeGe74oIIAjLjFV
p6hVbW3DWxY75Iag0MPKujEWZsOxL8LLs7tn1tQoqX+NCyzUNYrxvS58eC1YQWnt
4rmy+45jWZNrZKmTvubpMW/a4rCOc8mqHJ3bBiMxMxepr+aRI9qXbcqkkeluvbI0
s8muu1wW5oyBEZ80Yzy9zHZCFY46P8q5f++wolXhyfMCM4mQnDzP7dFp2dzVetyi
4ewwanuxxVtBiZOyDGZcYBR03rJWZL1drtsUVJqqddzkjFjqQQoAPMvLXg/2aKss
y/uWQlAz2ZkRmf9946rFH/XDHyx+pya+tm1IcyDEnOpb2kGG7HUKjepjroxuUyop
AcXSURmPHXrocrKwpgKFNT/aQVxvHmoOx4hAO28OYCjQdHDJNO+WzsAVVGZLh+o/
g56BkXQYxHFU7FYCN0tfAy4FOD3ridkU70nl13/UPIHeZvLmXMjExA3viSv6vPnK
NOKHcdKwb70XDOtcxJZf8cl5KZWu7szl7e3kAVjcA2XCWgxPDhaO1MZnIGSnWVoZ
pQLzHFcbHbPoQl55mr37AE976+5s6CZYaBCm8P/vkwnSYlUbZXQKN0xP0KnxpZXv
lsmFxeCVnxZEzVMnM+Z8VKkdm+/n1EEayeylYh1ICQobdUnHp5M+Ui1q/xg2Pbwp
2Vcxaffhoc6LF+AR10zeN9ZRoQ9kLdCOgE7a6p4C4MK7EmhJnYQYbftm90EWlnnB
WpDBhjRxSgTBgFOQTqx4TUaXUGQVGvH/AniqQ2uIORQ4SeY2rMpEDC9K03htMBB/
YYkSaH9GQet3dhoxjybeb9mnzH3qCBgVvOfskVFwTLhUBJ1UnrLQ/XitcImSq+m4
S7XpDTm0RwIdpWgVQbMRtH/mdC1B+lMLUCFRl5RGDGbeAW3z3a72hpPmezq/eHmW
n/qV5jfeQPWfM63u6XxfSB5pWKfHaKo9XjJDmFyDmg9TroJr6x7HplFofVINpAJk
xbkBDju8T2fP7nz9eX+9OGQ4ALfIEwe/X2NB3UbRHAescFjSVuHnkCpYveZJS665
9XCQuo1ttEX4Jkn7MGxSjnp0EtbWNwWoEiqznafdlR9DX3Tn7YHbeniqEI3NErwC
1F7gS/giOmWtHrCIr0Ewxl/OdnMxFlXggWdU41YxKb7jyF28eHWV3nfUV0xoDdRB
Xn3BIByU4vCBraXcN72TOTUxBjINP80ioLEJpMO6sLASLOhkrUs3Y80O5u04n9GK
m2S2va13E9oMmpfd+FRz7wY2cK+Ry66UtsmNbc6ac4FVILkEyeIi94Z2iMVxswqW
ucRyI3Xufi9XpS9nwX0Tr4IYG8yaD5M0GY5gFctEi9nkwNP573iK1rLfs6wqcudT
PG/kYPUt14US+vpq4Yt82oNL66EJr+pA554m4VIbC8z3ypfhi9iF08qABDAnd82r
sOs552sm5S1WNvJxHPu/VTk5FujUkZYIbXQOeTDXNcylJI+x7e2F4rnGBT0CMmY7
DgaVkVodId+u+fM6DBLSari4FBueh8IVTH9H0f6Dj3iIB9tAW2wqDX7QYEhrU5WS
HVmk3/gp5LnD4Lc99iNAXIefwvMoeui+cBHndhpYxrAk3i47Xz1YXiQqoFuD6NFq
uBBGQ11g2RyS06VU8/l/fRZFPlVpDfIFXApRLXhCn3n0wDVPC+w524TYkwlTvNIV
xJ+4044+xT1vjqrBEUNUejgTm1YGco9z07QxeAonutU4jlrpxBjDbu0u8HsLhmPT
q5KcI+YXym756DtuVEoYk30qNFRp1/HUD+FLqXJzCk2sEZnCKSREGDdmwlgDj12P
Pc13MC9BYXX0qEJM0qd4PM6bi/N3GHEcJkEYmLz847EmbA3F+bMTt+CN9dZOYuLu
Mqjq21iAizeFPbJ2SUXsjEL11jYiL3qRDvvfYj/frCe0IlyvFEhoGXQzwDPEseoU
JRAMpbL4JPvqP46vvk6soio8+3984ZpSOzqdOcMLVeskiNxyHUo5/ihRzadLClcU
7AegRMfPEN6z44Z0lrqZK6MAXDqKOqQHKsZyGvpKoktUcnz55lfbsbsM39HjZ16W
X9vQEpt+kc3HOa+RU575WE8G03/F8tjttV60DmfBCOuwVKp2NSRlQDbE34CmZ2vj
MaIkYjRU+WSXUq1JDbMAwJWzJhixyPXd2ps09jHGkTVbUzeSu66xIOvhUNi9CIFv
ZSzyPNxrFnN+B3NKqTD0LW1EhKlpijoaH32Mh1LmDNZ/K8w9hq+OzfmZriFnJtg+
tuasgVhm8TEn8Nbg6OYyzPhWtK0jSiVazik2RtpIVPnLwcZBcw0h4tv9MqSXKr5m
OawsfXYUgQSSn8yYRUwsd7V/uBj3XTk/ZdYxpvNE+1BmBl6FgBrriluxOL1HHekU
MKz+OiwCnCEWyKTm5CSlh4ZmbsuMK1lDJkg0ZkhuUto+1UxCv+glDsjxxTTBsC54
UvpOPU3GC1eL/+TF2zNNZfA/4hDtXs+J6FQROjGpnrUlj+C2/bGN9qMQbvl0IYyE
4YJ4emJHDO2bUrnLEfDP7lTb8OS7Xn46Ww0sBw1wSKcUmIzebQjTraHDBBwfvrqP
Zb45wa6zXJi3WaZWsxZi3AGYdz8CFLK2LM17lo3me1F6BFr22Bg6V0Oe3gvDxxlK
jbvlldfdBDiDee5MfLVd1MfKQ6xZc+Qdj+JX79oa55WHKHAiywURSXFUn3FZ3ugk
3NgEOAr0XKNRbfURJ7AKaH5dQ4lzNWEGKHcuOo6mErj0DAznWDSyiWWUgQ7Ry3iJ
sQlMfyiT67gMux3pBsnLgpJ50Vpb1Z9y5ly6q+YDwoxEoL73mP9uHJgxKT0o7POo
WfWtv/A33MtzEbFSwq5gqc6bVsrYqhG/vUA5C2FmYliZs2qDOzKwTmXcKZO/b+g8
GiRfqDwMzqcXupOiqy7z9gZdY9HNjUBFTfJUbBmy9hRtVeR8BI6zk41ZB+z2oSh2
0LN//7AbS/r0S4mAWrGNS3ASBSHR54B8aFR2/twCvbfDVGVanSnH5KWFTgC3HyTR
WqpEd1Tx5c56S2hKhHhSHrmy1BtV7ATAiYuHjkACNUfgJvWvH+iMzPF91JBe/4U+
wnt27t95V+J1NNt0h1S56JYPIfjsWj8BRDUD1LloCGzlttH2Vlcm7tnt4OE/PfLh
n4vPuDbjCqJEmYsrPOdNAUiVcixZDO3Cpk4u5lHx/vZ0d89Lt3FEXzQQ36igZFpw
eIVYI4HodpNwC1uIUFoefZce2y8HwcQdsf5ansi7VWdACWv7VrIGlNUPHBCQmKLp
O5tSXOHLFLotkpeXbfs7c6xa2WhjhLnaCD8zYuisyylDF3e5qcCS/0RLEbTcyoEH
SZG60TRKK+v7e619fg2BFsXg5jZ+ZGM1XfDg3gcffsEfFJJp37mMmhi1FcU+2pXU
wkwRoZ2Kv+bgg3+ER35oaohQ5QdlOz4dRfqvArh5r5mmnA1nPbTJ62hYCYS+SlJt
DhEC5DXndBAETGvGgl6fMM98UJ2n6TY6JEOoRgXZxZPaeDTMii0RW3VboDwEuYB7
jdVh+M5cLQzIzSEEeEOvA0/m1Ie/vaWzLHEWjtz7aSD9zcEcy4OuLz4QPeRAZNsO
DEBNuIqAyXszAKtqPH7SLeFoYTfuIPkqRWD13sZ2BEc2m+WQbzJ42H5sTzwSAMsA
1WNtUUPScjIRm128Cw5dMLzKAJLU3tCRLJhTx2U4pE7QIblLb5PaEvHVu24SZBsp
Myp+LU7zK+AlI8uI6Y7hAIDi9+a1A9/4hoJra+Lhi8tI1YAndw21i3IiUN7oZgDA
o0ecyJdSFzYRSZoEY0VFEIgyosCdvCMVh2hgIjP2La08F21cxZUkIwUqf/ovjDNy
euO5GTNw5HmAEp+Sux/g5Jhk8n0vs990XRPCB964xTdjXc3jfDcI7EUqFdJzIJ9v
JjjM69GZrj4KQc3NOpsSsLa1aKWA9lEyLcJjl2HVz999QxlmaaLsh+1htOSjUTrO
GadpuAFZfv2CYJJQqUip+aF9dut0m1jzIjsJQQjfnZLToE/lZpYW5N+SflntqfDI
aUzU4xgaM2j04ZQ/+44LLCqJBye/iaEKaq7nOMYsBusCTGs36seGuW05y4V5q5RD
jg+MguKPMEiB4uwoxSOyEYSpFCmUXwllJ19tvBv8RVtDXeCXJt3LGqcjItg3c5UO
utGMSqUSVJCCIOzDOUyGZzIyQ+Ifi7548+NiqvOLF9WdQp6HeWod/OFMs6IILTvW
PqmXtkS6ScvM2X1Athp1jC9AsSCjhcOpitFOO5p9ZuGgqvNKh+MK5COHnow5pgyz
XtrmCKpSTq9yOiAJ6kdkMh7xS8pzFQ8TlJ2vPigAbiGngqdJ4mwc1KY2BsXlJz/o
4gQqpBnaSyrNdjeGTsWAUJmQupQRYgN7otsDYNyjZ9oFXSyHCNNZ53415lgGJh7K
CHoSNTLgRuEpnCYWZUFe7kgD2eE6Fyak7RsgPGqkne6ZXFVOfzdDlpvdP9IjzQNO
ib+PrGHkmXT2GLxSMIhQpGQS7i98XGlrSxwK7urUvaT+3ri1O5VUVcOmr+DMvw9D
JuGpC7oCMpw8UOZD8AdVdwu1XTZrtRMifvZOKu5aWhye3LRT+YQLkndxe7kl2bdl
P98Uo5lx0JzpHCUXnAGBggKa1V3f7OGSeWcNN8ONQOks9l7oDnCfulrFQN7g8aD3
y4TflNUAe6AFI7rpJXdlw6k3LGJohzq7hTzewsHAjP4vflqv2+rDjhtCTZnKhgob
ryOyaZhofLTpHpZj7HeDVK1XaFd7pjGZZYTq54JfqCMJG7Hh5Vif4KW1QbG7k/QT
C4QpTq0lR+Qx04W4yM/6+47DJL2V2cC4CpifHFddJuQzPzsuorkqABV/nRcrj1qQ
u/L9tu3dHmZ7vu69kXddHElGvrNNiONCJLsaFe6KEo2eGRF3LtRVnzKbFkoJrhtZ
5UtSrdheRECTTeViTMqE4XQoXOyl+7te3hkwatAY1F7WQQ5xbmk+HO+MqbOcOtik
g/trwoTQJbUlgxweH9GR/3XVlPRaR5gy8Zb7RiG4xWhAx/O28xswVGm/ktpqddGM
CMWuecFGl55pljV7YNAyHT2xF60RfCHGZjH8nV/ZlG3tEyNEE7HVlVG9ikT0U8oM
aFDdFScPBjZYeCtmy+SOAk//PGPp888o2le2vxZ2S5d2Os5pgQT+w6JC5u4GIzvU
ZufUnzmeJlGf0YOoa9182OsmdbwBCKtpOmJR/jxjrHICOspxSCLGiT2qfv84TdS2
y3H7RccTBo15Rq2C/wQd4i3PFk8xIkWRFR0H2fet2vhWAzgyNTl3Qg7ddqyQVQie
wNBxrI4TuJ47q9oQrnYQn4k80zWJBfR6gQIr7F3wRbstx4oJ6ZFMswY73nvqjJKG
N2/0qPpmLvaTDspQPUMqF6rYx8+Jxri4AO17/eKohzUfVJWUlupnl+IN6/7MFMr+
DrppjrtivHJ9rdLQfW2uifuysrJjWSgwX8hX8wi0fqMOmwsZ9TRZn36IRWn/RMn0
H65XXYaj9NUlnWMzQuRfsahGUf0sLsZ9lSrJOg9UxWaMcJgCu40bD1aNAl4KB1I9
cdUWIn0flIfOhztRjgv/AzmbT4ebzAD5WfYF0E8CHQ2lDqFFbZUbCU9TMgnIE6k+
1Y7u3zzGqZiFogpRlpBkNEADwv1rBHlfnMRpysQR2cqBFKdsN+8MAfkJjIspZ5/w
j+OyVqeCF9XOugMCN21eJgweTNNCsnnx+tpYYoDYhLY5ez/G8ZoysMjUEODJgf4B
QOqWjkLiTmk8TyaLSUzQKwkc/A/nX4NSk+dABVRt9ZS00Hnd10ZnYNUViWwKpaPH
1r0dBZJeWi3ePonrqqLihZE7NgiNz704jiFOb0Oe4H6UFalRrRcMuJfasxEA6dm6
Td2nqXN2wYkD1MWP6F9h8e6pwtc2dg5Yt2K4IgDi5TFpBuGoYefUBD/Uhc6OuQ+8
RfL33j1mNtwsZVMoHxZRKzcDNhd1Juaj9hszxIX7FtcusJh9w1DgmXKASd/glAPG
Lhxxcu6iNwxQryX0SvGK3ctKhoQVyLyvCXmrdK8mGSy7RtwzqmssdwOnBEgLwkjH
rvEaPcGt8Qp2vzSUkkI7TZHoyd93PWA9Lbw+yPJtJHSEZJyI+0KRVEb+VLZSZuyi
Lo11U2RIVZJvMdYStDwJwOEZgRmbgCJmB7SakdQACj8P9BgtQBbwIhi+dFerjz/o
XQJCY4nllx94xrm8DKsNQcucFRz0/Asf8NlFddkvLGK+I2bKKsCc0KMQ/xPgrAYN
y8aoBU0JpMzYXQBVSBizGL57PoJMqZ2Ncgr0J0k/ghcHanRuO5Ju7GIoGxAL8KpJ
+fevWOhO0Fa4jW/EVlefEHgyZGv9Fk0lOHKx4pevgNeY+Lk5BNUt+xYKc3XBYMW3
9z47sUxovEfJ005UA/xZRO70OUECwZR0ybSYZ/13NJFliL+EmVvm4ubJGSM7NZGq
MWaQEIo/frTKBLbW9rpVhe9WrI9+sK857PqIkRYprCWDFRx3wUvmsWvgqPU4vCwJ
MyeakVCMThsYM31UMxfz+2erfb7azoZqovsdc7JodTnjlUiHaD4iaD3DAn0q/a44
xZAIVn1OurLSpSr/7TVvh+a4fDGQkd2NZkLEvSt78AnPfHdLyWZhXBc85XOaU8WD
4lq3j1l4LLm199AIXGqCHS6GkS9WcZKOU4Q7IZEW6067j33TJlICyaBd/AIoFNHg
nzvvZ4KzJpLpYLAYHW//Gps5rSNZjWpzkDQ/9mVu3+qiXww5NeFc/7J6VOf5DO2X
dPpksoIqi5fSuIWM9j7ACAj4FRTflWHlEfRNhDHbLOOq/fAqhyiMiS6hWs/Ml22Z
Sllph3xBksXnxNrpdZumnByMGfHs31URkP6O36Ogf3o+xn77d5Qy8agPzQhRwFw+
KBGko2vxbuj/8ZbHVJSIuUBOUVw1pjCnru18ZisZ40CeqOKvYurHmPJbHe1DoNtG
GvKWQNSNN8aX503DrWQxuaGgZmaGIqco8vY9FuIl4JZctkKuhmf3kqCbAAv6LinS
fbx/J5iaQ/rsecK4qFi5qjIkIVW9v2SQWEEjAuaKTlrYoaIizDWFuK45XhRf35EY
Lt/5ZMyVwMtDeeNCvkCadynQFhXCEhtcuTvyWT7yQVMzltIvxyFe7swtqNfUppx1
ZpNdeUBACS42rC7J2ehL7zYAT5UPWMbJWRMV5l02XoCNOCn4F39T24SAPP+yc1Fv
fxRkzerBje+0iq/6StXLi2nZRRSHyaZR2Hg8doDC3ZFmvNYUTt5dzYQzohh27Qih
5rrHQyQcyxGUa1p8Ilym6F1zDv5C8gLX/Ffg9xlLPF7kdlUqEW/ye7vAK8FBxbAz
OpPybwHRmXFj0JQa74uOENAMXIw6iKyP2oQFVWTJ5sKjHUogIUogHH3Jsw4MLfoX
MGGxRU2TRSQNJZkwoTj6U4MPslEyCucNEgUuxPAEUyOGAaYU6cdhnJ4SS5FuzDj0
0qlUwjSNLhK8s05FiHOpDBt6EnKg7kRnKSpXaDEukP21npFFdqr6O8LA3qYJYdL4
Yy67DEEVcGbL8anm3udTNjdMCeF+GHESsG2eYASUYwWbqZRYhp9fpCerOzJO74vX
ilTyemAaylU+o4T7yS5FWuQLebGHYNFUEvSyTpnRWKYMbK8vwB7331dno8m9rtd5
/qDH+wJQbKAJ36idQ/wuDp2P7BHWtFPcQQi+ivy+Vccf2NSAUMedkJ4UqXXz0PVH
OERch+OSaVHXMKm3bjIk8nWsvyKP0qGM4mg9/0oG2KPOdYLK8wKIylRI/vIRYW0u
H5Tnww5B/6yvvZMecQZZSKbw+z6GmVWwQFz3Skjbfow2kgJUiozNQ9N2KIgz/v4P
8S7gZ5mAeW5rxe6n+s1V3k4VsWxiuiYZg5QfuIPE3vghfI0dXDJd5M4dxyiuM+y0
AXbOhS8Qo9FHqJBzmGwMTB2EDWw1kIAJuS9YpvoMxh09yqYKFd5mGQCEph60h8XO
K4M0t00Bh+GzHLPH0zsuib+xrq0pvTLSQS9beMb++s9F8jWsLjwH9MlweKSzxL0r
rXtsYmd7gAnFPpevJb014cCQdu+24IzjAEScRbtfrARZyLfog50cFMgjsJnmfLZM
vX4PEUPM/yZNT4QapNBaEoT5+8GLr4flgfpqAxKmVkEqZivUvy0ow4LKTR0C6pgi
6756+ICYya6DuJAJyVNiCXXNAbtwYjUCOfv/I4X6w8xblX6n7K7uVS2re2xHoi//
/uEVdtogvTW7/4lXRSXyDzTEy8WDplzMm19zSULVYrFRu19upAxZQjSEwqp9PeIM
j2EsInnoJcsDLPAkn9XM+B/4RG9z0Z6wMO06NQmPn823nTAKWrYoRLKnwQeQtcy1
4TWCXVi4+Y9nqcIunzw3qgGYa3MKSkGOQZSkMKPjJb5CjUCmgveLpcABPfIJj1UY
itiMBl6Y8HNWhBJEcjfAosUIft0C3ssyS09iXy9vPXbfVYvDLmnZRhe3XF8Skgym
GeS5GzaXFpfgwTNBLyDg49eOQWnfH23V5jWDtNSOVZ+i+Wf5QqkwVOBRoti3z0oK
vnljQ4iDIe/YxlHfrOsTMPcQtYFsyKlO3i4GxpTTGW33QHKS4blP74+tTwrT7fOh
U6waBxCkHtKb1LsL3ruPoFdG0CpI6yAWEQGDfdJm6x/OcvPC3ThrUasrRYzfJEFW
HkcXgivjR6w6f4vBTvBI+FCf/9TfPcTLdROh/SJo2Evdnae03Ol8lvs7K7TurNbB
flUwLpYQDv5dcCU5Wv5hzkoPDvVnsMCezdCnZ3FpnN1wY7LniEF5MCWTjss2KG0N
Q3OEorIbLe7bwmfpff5eG8FhCubD07IeIe4KC5hdWhC/GRxQRl8M2VIMMpRHfOZ9
1OLbgBvpELc/Hc4XNGx9vYaO0z9OPsIlvohtHSfJewLmKZt+ghp+2odKwA3vwYMw
/ect4Ljrlupkel1K+DyXHsaSCSwujB//Cvx4yr56UlmTx4iqVrpSIcEi4MeyBmBK
1wK7xlJx/8xrKPWSZD6+4RoE/I5tnhk1cwM4eqS20eGu7zSlkiSD7yytv/pP+Em8
fK1AJ4wlUc/Cu8FAe1ELH775+5LoHlwQTdK79X7AU36oyld+D3JpNsCEBG6paXSj
+JofavSS73Ihagro45s6KzABlekFgN5+55awfRPh9i/5RJz7ETatyq2nTob6I1hX
T3+TJ9BTcLlj2/DGGMDoMviTNYqHDxoDycvjrD6b44U7f7Ws2JwbBYOTLiMfgO2u
9p+koTymOo9EAF4BCsr6QVUqfhFHYMks2vsgPCxNK7je7I0CP8ibLFqynRTmX4FN
8aNJEIUeAdc/Qc/Syb473ilj8+VHZGiAy/fURC95fvvXuTCY2uUc8bZSqOX7Nb0H
SVycLFjDYiNlAlmJjbFYVZYMkJbsvLRieoX0ngnyG04TKgU0sINiVB4QIUwjtBCB
/dBTXLL/uy1CSDFPQm+BX0a8DMamyZyHIye/FNFxIzWqiirRg+wlZVWSHT+6RTjx
Bv1L2Ip/g/X7kmVKNK2zrZza7IP+lyjEoX3Wgeel6zu1C5a4CZMbZO6uvpUZtbzQ
SH4n11BTyz/zI+vm3j3g825VwFN8+zEvHAXYpHfZSHf/G18CT0uzdAC0xPeAWRxe
UulUTty89OKk/EBQyp8ujOBkY9jcOGFqiRXfi2nRs0IlmFxiaBYKTlNXnx4/Kogi
uZgA181amL7lyZApmfrI6U0UPcVvdh+zkMB27hK4FioBzo1MwB0WGGEugG+wyjRo
6Gcgw4k9INasaqWRHvId3MCJ678snMk5ef2lC2dLgkTbSMW4yCZMM21fWUpW4roN
YeAJM1+UZP60GAvzd9ADUSFV9SoXw+wY9FyZyReNUpIgOkrIFYgpDKzmTgcaw4Qj
3PumcwJ0cDaD+R6uRYPAiNtbRcmQT5dMluTHvQgIPJPebhlxQmQZOApg34I2i/Oi
d50qG2PJcFIT26MHIbUeVlHnFYvPfQCmi1d1JsTnvqWX13BTDYo3FevipuUolpp7
ySSqyGFyCnroHFS9J3LokoXn+Q6tkwowFCEftqf1hULmC0zxZQH3/bkHQ0yzx5Yg
FUKP85t5njw1P22mXpHVkA32DaQUQZnBROjI2CPZrfOXl2tbJfLQlKUPPunq7tz+
+iOZUh2Uvfka89303JBLwVUAulsWqM7kyOgKgkqro15kKUoZsgdOavbR4HtJ5tnX
GVHCGAb91L8DAdDqj/HHictd7yvG/Hbi+qsRoEouTSFnRFrn/9x/a9QK4ii4H6iB
K7rzvdbnJE4+gHZnBy+U1GA2o10w1lehVuaR2/SYp4FixT3KveTW8PVziCm1qCKv
/LniMUXM9TIqOYT5Z5OiEv23GyXzHLYnrYnJgc4SDE5rkbRA4ooFX1fUIjz3jEys
TEmW0FCpkGsJDWfV/64DUQJ/jdKwNdJ8jowZ+HnQ+kxD621BS+HVmbjUi+Q6/VU+
LlmBpffWzHr5DHn3G8bDfoOlUppM90ysbR7GEvHaQ8X/n16CIMl60C5aKkH658g7
iyBVdWcAKS69Z9rGcVXahxYe4Rgaa6zdV0EKiwxJpiqe7N1O/HKHM3NtdlAo8X19
KYdJ0I6sTqyJv73IwhjnmDES3Dm8PyHbzJrk/kjk6TN6sm8JB7SZPQ1+jKIBTzeC
EtSun15y91zEL6R9SO2WzZe/TLIFbVh0TLA07OWznvVbDgpDrcLej5u+v9DZzfjP
7LVu2z1UDMCRbQUD+J9VjjVmXJzgseb2PUAiZcpRQxNEWQ4upqyrLijnWHdrlV+f
uMJz9JHo2LefNHs9aYGn2yboRjG2Ml/uAg7azsm9LSrDw/KKGBfXq3KEP8NdaO7K
c0a/kojzTmQNPgaJ1m0yNGqoYGhSj6wNEcu1K+VMKGvaLvyjHznrUnZ2LKbiUDN8
3nfTbk3vqW00Gawonxyidpb2vpENU0UDJwBxteQ0kxWezSYd3bIrEGGo8/wd/ohV
uVdjdlJnii/CgRH+cxxCLghavUYwziObBEh+BjzIKMlsoTr3H12F/6A4xPeEsdGb
1jLSyquGQVI8vRPAMUebHRWFg4bdHBntK4YTvk6oaohWIw7/HO/sVryywh419KCY
gB84P61jjHwXg70RAX7M+2nmVaVj6YJKf3rXZu10albySy2VCc1tA7jXTC9pGEJx
VIS+WAghrsh7dzy2Udj4qjjxXqZkaUPGnPQ7e77LmJcXOHmasQIVA+B+Ia3ZijjQ
SVsEZU+NzGfdarVaCNqk/TWxWwgH3IojpR+ZgPPmMCsKtssOeG9chy1GCOWy6wMc
q+0/qWwGF6N3xMBdIywtNZE1PubhKRLqU5Kq0YwNc1TXjBatKSwrU+mk92UGSXk5
qBWcJj40folf6txuTyx/YUsUcyHBzW0zKAJRA6b7nE4/SwUAbVgJzrOnnKpyPL0Q
FNqnYHa0EACuYTtUjbK+mwrQJoL31YrCNc5peRLnJ7uWKhBXNYVumKkiPdf2nEOp
zlqRw9hHyarxv6wblrcGZue5UUTybLB1UAkhheczt6oe8slAzF5zeyYkyxf5nA5u
/V4JFtubxNEfvKlxxO83T97cA3qeA2WNSBY4CYL1mfYuHf6n3xRGMbFcfy+lKQUF
7NgaKXr2mUTOBULKM6kXBH77cdJjTXSPna2tnjqs3IpRQWR7OliIgHCNYQt3vcMP
0mXlNsMwjTdJFC+OYanm6WIjGUFP1Q4Q7pZw4U0CLPcEmI2hfUy1dH5s9m/n+Ib1
gyUyn9pSHsz18H3i8IDtoqTxTxngoE0WapCMZ3jCbES8dcV3QNqnAYIrMThPnGGf
6EozgwGV2gg9Bn/lEE7CoDpAHScXOhxJn9QF80TrhTIq0HMN7pz1GAXdkhqjvgVl
Ld1v9Xif15NUOtf0tzLX6eie04QevvadiftC8PPnI+iKn83nNj9CfzBOodEzK2tR
yqIU6Lp57isXu6ip0vmL0V2hQkbVmzCnY3Yz/3BCs7QP8NopCHHxrmuRDtX1rg6R
VjxcCnqVQ90IfuBItJ3r7aKSIYQNVDMbXPbjcaZs01vmXRqCerOmekBFo2SBGi0L
E3qvSYvVs67B6M/cxvIV3QthYrFzAt7eaymn46mYH99pDPM7m6FxNYJqWIxpa9ik
m0AQOOlfnmOESEW39BzItG1A9fmtI/T3UkQ0EEKBj6apiW+IP0Fe+bJznvbG8FbF
EIXOyh4AE7c/erim3uW6nPChLnFZuU5Gj5PUF8ldCcBg7o7B9v7BTDhuMF6VAtiv
cw5voBhfnuPxGN7CZVuFebv/AEJQJx3Kb/L88+o6O/tzaSlI8Rpy+coVU3+V5C//
ectNzmT4Lr2CKoT363wXbxKiK4ZuoTRBrU63+iJUWKnPgRvZwwws58ealyA7Bs+q
GZzBe2qkXPQkFqq7aZcsE4l8H/Q1KM3cSB+ktED4yguXE8StAmtXBW2d22uOIqeV
F8JkzxqkyYqc6XzO9jXP5C29nbGike4vl0dwUCAs66Hbiw1u+inJteTarkm1dsqK
xTIjA9LylKvLrlzvrpXAwfEPmxQ5Jam4ZYysu111s5senZpmD5mxJTBTkaHZ2/LV
iVZ8rWMcjZtzqrI3f1PKDHbm3F0vD9KrTqL3Fq4K3l1xfbb35Q+Sqb+hPo8Mibg6
VGCKNXtG3uJVjIKR7jPu6gZ+iU2tQFhCkSQanBJ+eofwY9FHYDSRnfRBiIT6KtxT
IxEXikBx6HZBNJxsPfE8lnO5sn1s6AyJHV8jaYsM1YHdbAPo42iwrYTCDFFdZUPG
NcU9IPdODPOwZvo9NdlwgKbTWijueokAP5AnjG4ucvLtTBqcB/aM5IBnfYxLJq1C
Q9KRK1AwU1L3FrmZ/p7LKwQfd3H5k1hfT+BDjGmouksEud63eq5iV+QmWwoGC8aO
ws9SZa1lNXYm/9qomxBFJIXax4j6TMWK6xFBiSS0nHVakiB/bjrKiOf3FnS/nPx1
NBOp2Tp0B36fPOp70Ne0M2qaVYo1bZ8o4RhPbWmEKMVrVNVqDxYQwaljLUjPNuL+
C3MMRgI5KDUuWi2rP0LCHo3XVI6hbBrAZDXj4nx8sDluuPav1QG20tIoRqT2VaPs
m3pxquOuieN0b6M/glCKxoZteYbUxu/k4yq95UyMAWPHTmVprEl77SVHi2qpLO0A
Pk+ByKhViCHlx6An2G3ITG/mo8446zjJY50uD0EaeI3Ac3vLKc4rkzq/jZaFNkhI
7jMBKZBuBC5uT16arwY8SMNyQxRTHzpOEdHvcdOT8MHl2JSn8AA6MDBV365HGkmI
kUM/MiW/ElmW96hG7A4uEe+sEDTRt5Mk1Kcpp9NJJA+zCy33Vqa9upJwRv/G8kUa
q4lzEw1Pn/myNFVOoIz4q2Ej9YiwIL8J/7u9THK8+Nry4ictTbdUOKLOrQ4kvf3T
H/5/PEp2Qx1ZzhDtAY2UZ7lHhHpdqBNXdBbPOx/NfRiRxzHMX0+X9nFZ1G6NpeXa
xDWcGGOOslFvORN6031f6bdSW7WkzMbGExx2gCOywIn52xWuCUwUNJoCZL6BEt2C
kahgxetasziUeldKVLFx+kUkIywtdej15Ea3dcXLgBTri7JoDkSOSuTmvoREBq9J
vYSVRP8CM69nQReqX/zn4ahuEENdALqTZ/zdQMvpLpNJRukF6y6HiqjXK+39dk/u
56Z0thBqyPm7X+amyoWNMU8UlDHpJyIZEANnniqM1796D/rsKwPyBU9ePCGYuoxZ
kw4qIpaxbyeL3lPOzgfcwjA2NBIHVBSr9Ge3i8Foo51+3jyTb6ajOAhdt2+YHl6e
vlg4izwtaPuoSmevwCXSDFQB3U0+1Y8rjRrDzGQ9YYCT5vau9ssVAwPg+Tzaitzl
vrtlvd3sNgT8pCJ5FZkD0SsNsdvOQMPm9rttN454OmTZtQChPT1HbjhjPb/woR0K
ihO1pbzcSPlGR+MNDSKtBCmunh45toJpR33QkMVRrwZ6Yita//LGvyQZZoCwqjIx
9wGkMVJ3B20tFokF7kmy/pe/Xj6su9KezmfbnVw5tuNHGCGUeoKgvoTUs7KrB73W
aZHCXB174Cl2EzntR4vTkESXCR78dRT4MgCvLA3wPU+2nsCRvDUwIW2VYnGvMGFO
GjKqdhGlfjYpo0sqLPGqCUmTAHHoRc7KFOZrnNdqCHRX3v86CLCrS2oJu/pIhFeb
/mR7x7+Urp8wrZxxyqrgkbEQuDO5p9u0qhRHPOlr/02grSkaFsS+qFQ9Y8zRH1gw
q7kSGzE5d7zddwbeFsgORY99JTy2uwci/WMbMSeH8+ijJykzyP/xHsQ2ia7wzoZs
aPwNxvSDkmXgWbXfyMDSPkOsc6Op/l8xgFOivaWgEk9XWtyeENrY+Hp8R1oQBtUa
1ogQEIgV77yRK59Km72R2xcKdicGcnr00S7VSH61fU3oyHjTgxXiaYtJjDQYO8tF
VLM+IU4RAGb2/Nsb8VRnSMveGJvey8Ia1hXvUbFGU7LPdD2pzJG0Z8rZqvTzKAQY
sLHwqtMEt6ZMq6fUz27vMq6ztXAb8pm1fQ/viGBC4drHZH3Uqe1cX9kXNMFQmv57
AsZRpi+QHa6GEmqbrtLWOfE3IKCV35oiZvWnz81ITVksLLe8fH7twxlxTmy6iB7b
8jKiG6vddAfSLIIFENtMoez+VcOaSpWB0xBfHwG39Xb0w3X96MY8okygDK8jHTJP
3L3S3pIQtlGah/i/HknfDAegGGrlkRC19kJCgTIplU7HI4P8tryu+pZtx5jp+eIB
kyhqywxp8IycqesZgITZV+lVFaIo9KW8SKF92N0jPx4PW3Dnhhj1EKT8BdLyzyWD
CXzZPEEj/Q7kfGsL1hS7oz6OR8UdX3dkeDOcAe4cX+Fto7F7dRV9PFRVMwhBjNx6
RWONyAEhvK8lah4PICcrSEvfqrVbCAM0JAvFRDBS7wp1sXlYN6tTzT7i99xGr2UR
5GhaHVlutbQdPvdK4eal/ngk8rZ6zZT6cwXuDpbHNjw5FyOnFuFUP+3SBGQJnW7H
YXyjBS5pM560gFlL5LSlvSLnZmCL8J/txFsPpoHLpWOAnPPeekFzID7/KhAx9H70
Wo4f9AaG839zR6MHR/wAX4s/GOGVUsl6YIigYdnMus0WKck56PLKlgXhp4m4hCsl
IPlLldvLRY6jtrV7645kao2T8p1pW4nkkKZZXNgjSD/RvLw8zgRCEnSDcJ2AgtzJ
ckqVlDf/aGzLLNPZV2REjfaSKe9PSn33A9h06V2mMARKq+RPHKp2NYVlui0la5+W
gzZmPhGTmwA9bMO2gCUpsdq0J5/DyEdB+GJj2pOn6S1PruxygSXw3FlaZICrSAtH
HKqRRspIrsyfd89oAjudX46dQliypVA9gTHi+JuR3feu4hslzZI89T/80BJ+txFm
mIid2s+8LafHiH8dtp8jE05NoSa6I2YbmrKG+AEuiV+Lm6LXT7Xn3PvCwP4/8b5g
XY7Xy7XftYWnwwg1VZzzailGVKOEtLj1cDZqUNlF6FBNuwULVNLYBQx7BwpZc1ic
1ISmVxfD6xCwdu71TRkEUWakq2dUPNAfknZeLkp1cIwQlO3fHkB2X4Ar/99g4RfE
21TsquFphokvOwMLxeghRhTWZo2ty8l5lBsYI/UvPFzKJJcCNTi+Onu9BkY9abaf
1oUyq5Jiv7WfNEQ8eaJE+fpuvdPC6extMHySSn6o7gv+5dinoupn6j7yC5ZKLl4s
ysVgoXcjWd9CsKgBQpnSDP3JHn/i8RbMnF59EJbcc6XZ5C+Fs+zrpmSjP73l04Ek
+znjxustL9jpCHCIWbDiBuewesmPZlL2uIR7k/ZFJ7uDMMA5jQl2Qqozx3MF+awM
/ujvJjWtM0roWJDqxqZhp4sMrHSQX/4zCD9kQtDJKMCqTKLPZHuIVdi3c5/9voJp
xE9kpfwRw0Cj6LG09DhITgg7iQfbNOWpvPfZttVlUdyKCcuig189aGg0uiTFo/Qk
baf9k23oJdJVjZJCTZjSueOTVyP1WJ05Baer+K8a2UP6zy7/1KheLwVwwAWk6wYs
ms24LZpNwLqqCp2xzuHiyGpQO6F4RCoS5emRHsPrBHzNZQSLhUFG0KmzwPW/4JAb
OKQFuJQcV6a/ZG0uk049/5tkKrJ4VxIZHlUArllyfAgpJ0J+3cbOZ3i0Q+MTzxct
DUHwSUhVre/h6wp6XH4n8/rk7wroQDhRd3Gbwxc0i1lG1qnHri+to+CR3McQKo0X
8COPmGfkiqP/IH9/lAoY21UiPUdwPRkiC8LI1qrj/RQ7i/K6IS7cv7nFYEFhRGa2
EA5OmN6nEklKYEq2/f47i4y/3XfhvyH4r7j8VNBZDwAd39pR86+rRCxe+DCqJHDx
/uDXx49If46RC/QP6RbBwfdx/pOkBmmWTO7H0Somag5fYR2/IjbtGljR15z8zgok
p8tbHJS+6bkjh6qz18/A4AJyr5o5Wi0EzRoOacBI/FjVQIEdu/TTn0ycsiSXetw+
PtS2Sz/5Fa2+W/fsigBgMLo+YyownLyyi2OqhfHa0JzqSXSY0WbdnR+r93efcgfi
vEOhhVCDKcTYuNGIhRw6fZU6a8ltO+qTr8CMqKMz7ZMom0oyZZuk16Z6A5uWEozi
wTMs+Aeg4JeeMIb94796QLeMaRTWULHL2DAbJrzUOYxU6S5sqvNJcTw2ksu87mDO
QOVD/hbLWN/GtJIamvTg6xLUgmzg2LWnGOKxenIQHJ+fzZ9k7EGYE5oW8CcxlaM5
nAV8odTyTPOMIDo8bpN/w3BijRDE0Js66CrS4LYg7tzwRntJ9t71di79LEJJNGVm
YNYuiS8UeXz7X1Wpj+gQ+bJuuVAnrV/pcFfnaj/Sf9HRda+k12vqj4tBdLIARoRk
vlWpQOxSW24XJxBpNjUVBkk/eL3yVXgRg94oQT+LoMQkCCRYadNoHfqr0cLjmxaD
LDPajC5d+KGPg6G5WfzSyzE/Za5RMsFN8ytr3TMPctfvyf8dLcIkB8pcSeMdd1il
atKm8swMZQkRqvqF9tn6gFjG3nJ/EjKGaDLt4mugvW1rSnvikFlEedUWdWzU9FKV
Xr2CZVH+OI6aEV3uQZOV6lSh/6i1f4fo01GtPJDgoxvaAuN8vFnl8k52eokRC9S+
0/tn777d/auQlH+Y0Kr5cXtc/tRdhvwi3lAg3v3R0cbf//Pjd/9UoVF1mErLjadq
DTQxT1chSqYe67o/PbQhy+QQAOtrHd4WUm34+bY1MhIQ9xhpRa6COIsxk4QVUIwx
lC3ir+sVHWEOW8DCd8b7bVXg0YdjO4hn5/Zs5iTC64Qf/LjjJL1P0YQqErELGxYK
NiALdcuq/rcMz5AJt197wanS/1wTpvB6FKEHStTGxtqHUAtynwOrgKr4wFbMQg4O
T3OTFWG+2qHu5tjtS3ud8JmvLH5mk3B/vK5y4+PKdcrMMRmJuNZXpJQfDFVg0YUI
fTfkc9NmmX/65Czik3YXMLZlmUh7Yk/6YLhzz+4GU+XkR4rQoCZkBXDX75ufLx9L
Kl9xd6fTkLrBxJAbeMo92VqYdB3JWvnVaW2sXeLijRbnJkGgN0e+BVu08O/xWyhh
IU0jlhyyRI7PDSkR9mWo3g2TlZ04fP0NmlwznYpzqrm3+uRomRf1CVezRM2uXLju
sJC3+QAHFlFq0JktDZOUP+a/RPZHQ/txmZCEUl0ijA6sUbwvn5cId//zjKcRJM3g
TyfOY+Gc0CNC08kiImYvDLqPzN+cpWBzQh7rZVaUQXRaDKqHslTdcv9+sig7dxi0
Z8CHuk+XNs9nyMjxQgDPpd5DmI4i9ngHPwbGjF8DQtEADbgzAaf+mRr5JYsZUNmm
KVN1/bzGfjPBqs3I5VTvrbwcv0Zm61Nvx97Hmu9kjqCVvyQvpNABoCVYRi2OeZGr
INBZXi09e8U7GgdCaCsOJoywXTRGt2xSeZpWBcbDxVCjLrWJIENl5KDDd9CQp5Ld
vcSqH6hLjzwCV2gDE/g6yxa2Nyae5qyXUBa60kh2w1fefKkoFnAG9zOMuVhp7Dzu
B5HneIJnXdTpf5WsCMDNtXdazSFxBxLpQhlqUMqsYoncBH2AP/HfUa5sUYRAVK5l
IMIZORGTJ9b8POFJBemzjgw67A8Dy2dI/JiZiq7OAzg7fdPTDCMN4UyW9ZleLfKi
83XudjRU5cxIfDT4Ovz8WctZDzfATz8axINd3sCpitz8r9tl0SQeRuXCcOow8eVB
+Zdo1XARwuMoGPyj8HT6mXcGQVNVlzN0N+tYTzjxJ5GUqIKKBTzWktgUjCikfL7O
i06/9W6aWvqtGmTTvlU6mqBrxYEDEE1bb8zwN45t9fN16y0bSbcVUv66vtpFVYVE
Pn1Ko5Ue+nMBT8tOviVGuvA5S9Y1kzgja6KSpvPaRZcS5vbQYMp4b4QWCdTwqhL0
zN5j2sqB96haY7RF6SNJEbnfsYE4AJO6fqV052O8aS7iJJ5ys9cP4RsaeGFJV9Rd
j3HkxBhNS8LvasmcX0vLgxon1Io3ll3w7YhkMff30qsWuMsCcy7xZOXlfjbdFonc
Gy/8PbSTqlrrgXeHzdFNe/saRGQUQ0fahboEPPuPmG/FgBsZHZ2ACk01pXIk2FBw
YatBGme/ThpyPILIzhOXZtWWJv4zdjsSKdTqT+P+Ybh/Gu2SYYaIw9UjmjoSpU/U
ScWdXra2m0PjOE6JNdhkKDGTqtzYsE6gwk+yPFPL4NUoLHRkehsLhh572CSW6aY4
XcRCS+tnuzthBuiefKSUF1qfqCE7LSnyEa2NJl0x+qbeCP7CDhmIIHraYI2ppjpD
ZGCfvMvpxNQilk26Stok/rDPovAMnotyFUP+y0ssa5JOk7Snm9ecVHf0/uvIiK4T
cdHkRNZzALbVSbbru/0o8ogfIEPtte8T7CbLFonR4HUFjyXJ4JexAHRHJy65oEbi
poYo3bejmaWMdZEYXx9Skz3lZe1yAHeNFbeyB4f2WXCPx3oRn1WvM3N4MRDq6Bse
L9WOs1l75A51VkBsCPnHkT5cpP2ToFXjs4a9TowqeiGYn3ghHX0scsdEb3014kO6
7s0ER9PDl9enpZ74lmtskDaZjUj0x3ggzGOk8E+HpzDlFtkXoH5D6ZZcv+buddYD
2/vTOjWKJozqr6y11QHvgpjbLpmfE/Uc31XrJ/CnCyJHvu7bOT7oo6tfhcmYaQPp
LYsHgKOiWzew6qhvCjeYo4C7noVaMBjRqEh5IRlJgirIBmF5unamle3kmncM/oOb
iRtj7c9VQyV1BWeW1Zb6NXcZcdnLE/axeZSZ1HPXxodU3nrFzHpdWQ1/DGH8NDv3
9MywZ6wRNVL80gTTsgJb28TeiDMqgWsjCxcPZaw8jIQ2QmNY28aqiuRVCtKiWVDC
zvCyjBxYZROK0vBSaD+PS09ELNNb9eQHwkoldS7SFH1wzxzCAxl77Jn3608pdw2T
3sD4a2MusHZr//N43ACXQZWw65N8wdYmz3PViNpGYVHPaR4B2U7W4V1asppV36Dg
K6lBo9cnjMUXMOHa1wAqebkusLk0CaBAeDQ4LTebYYlTkpck/TZU+EwujDpMQh66
xagK2QKhmeQi5eEplGLSRPGcxai8jHZxRvzqe7MUaqBtZIKajh1XTMsUiCfAucgt
YPwwcqWORwApz1dKRbFsWSzr6VQjRn7MRor5CUdVlxNi6N/hhHiyDpAz07QvsqCo
tM2JZdTntE7JtkrFrI6JN6VjgDK4iPomdzEVF5mwL6dO/sOa3EuzkWJLCdm4dAiK
wSVXLh2vmoN5UH9LeZMRRT4fYfTKZah9SUpUhgEc2thpYq/ZyETPs5I6S83tyxGW
wQVWFmSjC3oFJXWN6Ivb16QNRJKDNJ0h+8XwA9kBiUgOi8beFUHcxBQJoViYjsij
QYoviDESoAk1ywfjb/9+hYL+vB4MWvJhyxNc2lrwySFZ7cxxwm4aJZtxGX/rtNUw
XVYusjSt2N9xcxTZGcIZfDeqUDXxAqWbYIcPBzqR2mHaOC52Q87nJg40URggGQw1
exPEIX72K4d6gEVG+WGolj9egcV8TxazHT/LU7ZLGNPPnUqqhEVgpgx32cbi1Gv3
0taibRBRkEAwVeX+tYiJfyzNtsdgkZKcExYoKkCiQZYB+39BRj394Pt4gTVfYUXu
Qej46bdIBB932H5DFARvnnafELrF4jhTsJ1zPGRJQapOrkZCWsB5fDQlboGPfDnE
xH0laYfzxDA2wqee5usltFbakV3GDmArJMv5HP89+ZNU5ym32T701aJuVVGm9xFY
9NfQ/Fj9qfp5s3vEsPQASJMKwk65li5cs39PyMRr2hfC5s+TfxP1UIW6qFW1mu4a
2eeDqefzciK2aYcJNLiDVso2cLjrRhtahCqYsJvoHIQR2orcBlZra8r69oVSw3Tw
geeK/cTXgYLZdYJ912k695/9CB5TiZkOUn80fzqjLrYqLliLXzmroPvjmRfBBl1K
Ak4M15gnZZQyF0bLtkDSTRYAnMrDZSSyEgKsjB3bm2xoLsnyC78rR13yqn9gDeSv
Sna4Oa+tonQI9T77MIzF49CcZQ1nMw04MvuY5yD6B0iHXCjxxjN8QgC1TzqRMIaL
t0wPn1ulm+vUHy+G4uZ4azyKVx+LG7Qf6YYFpf2nkCWWGgk5cAQTorV5ly93sbi8
fYuNEeFsfORmWO6paTGMGfkCgQSq8t5PyVzX5vOGDHz+VX2IQRZpd+iO1T96axmC
jXg5VnpSHdfIruL/sMkSd+2LAUrGTSyU2G5HIjCFnfV0zGSi0tQdCwCmocyENpKm
HrFuFFxTlzpwHYZkAz6Q2LxxkS1k+7aFHBfdB0MJWrigGnrZu4tX1ZWzg18gJ0un
b7+/6dhTv2QC6Pnvv08+NmNOGouZ7sh0i0DkvOAocXZ3r1BT41kvfC5Ydz9FV57M
TP70US3HDx2DfRKRwZ4zB9wXQb8XabRlBEpKalLUqPac/C9NO978TPzvFVWui0QV
Bh1xrLHKbhLDLOSVtqu1rMYXgsQVensL/X640Yu4p8pm+ejcvKBFywdp2iJMNSvA
ropj6250bdhQ2Zoq3EJGk1w/5XAho40R7RPsLwL6CZtvlLzK+OqsiZmdH0J02Vj4
HpvBbGe8zuYvDj7Y9NsQmb9KiMXXmUXDb/4kDAf+ohi0Hb9hnHc/TmPKz1aWpkkr
QC+Y5hJKDqDgBf9VbNzESbqlY0q7AELxWWoOYKcOCM0/Ol7Q09dyHt2aW61oswav
ZNYmf3tAqyKsEhnU2IkP1Ia6gLAXAvztP6rmOtr0Qrv/X7FY2lV/AHHqdcxGe4hg
biuBgxsSQcPYfNCsd2zzGbYAEpnRZU1omCR3bFN/7EiedHiumE25GeRSADENQtKZ
EeYbOjHJvWOioPg7p70u4pbi/BFXp9Z9humAR1VlgAb6wAre/xHIj4ZY5GSha2Y5
9cnutImlsMO6OChpwvEJv2bswwam2KCnyIwFhU/ZI87T5rE/8XwSHkH3WYqgve1i
/AEz33Tf44nObibLrbx+X1yc8xcxFQaDz3x5nE08TvRfORBaERpKLMZmeCICPLl+
07hgQ1LzoeWrPdbgEkJPUoZf3z5GFLR7kcs0WgReLewB25m/eXzWiPqh+2tDo2z7
Pl/hay19MHOTtNqubdryrDmhXVZfLix5glJ+RabsogSpDo9XuBwBvJzIxak7MdQi
EuoJGHeeL3GQYARow0E0OiiVVh9HPLqOQytvmvoTJTRWV8WWt8nj4jHaNAjMpb1V
kNyhTYqaEQiZuZ4A0bD2oyEbQVpc6VFO1+zfW3OcckkCeG2O7HYdWGWvTBDcUm2l
W6kxwwDvZy/S1S1nx+Bbh0Hwfe1x9JY9Ok+TnBoJgLuXPdDTjFI1u8Goq8SmYRiJ
IgXpOI0BP0akl82tFIbleYXH+dymZ9HnLgn04l9ngN/Bg3r6Idp1/x0VOxA1vLje
U+U32X1g7cgZ1y6SqUjUivKzt+61O3QJiyYlblTKDCqxNmrZjj5awDIxa7b/FFnk
EGOTgv0n6bF6yREMGI8eLCXBvYRomWQDXUHrWIkxBFThWq+eLEn994EbQyrBntwH
D0sN1hc3/KyyitCK6wpCwdtsFs0uJ8BoVyTmyay5E2dJIe3sGwcdGtEh0U7u8tB7
2JlFqILYxD7fHt7nWVGKel05N2KFTviOSA7RabipC5eiAN+hKSRpASW7TEzez4xq
aAB/C+P7Z+Xj5z/mFsF4mY8wv2PDoUN4+6pGsaxMOGASD69+tQnkOJoWEikHGQTo
Zk4nYr0CRiWou9sUYNj3Y17auWiUZdi2XBkqtWblka8skcbcjirZ1iatA7w9obKZ
+9Z8U+GWOUGOQayaxYfHVqvtkdYx4hsVWBNzVVMW24tjxeO0lyr6nuDQacVdLOTJ
z6O/aDZqTEpvtozWs46x6ocbDnerg5nDzbexfBSeq73ILz1lX5iZgXfbeh5OX15p
9m3RP8t/MJr2PsxxkyF8FZtPv8nJ1WhHQHhofZu/6ZkYiv3ykgKNsGOf/ys7D0vH
5lzXMQkkDdxkREdmE0S1+VUAFM0eMxAKX9tGIlJj+v0Ij1ZThLhAfC5RuAxKjTYR
FfLOIU0DXamrWGtBy3U/HyfXrl4z+L//wq2HXV2Q6r+R0WAOI5BH9D0RmiV1MVHh
04aINHYdygrb1wc8PvZpl4uEkCy+gf8t/CNm5TtOhY+T2ZxPMYrLpyfyMFO9YyRv
6ywHa0yq/abGyP4m8+LcWGDWz7/insosStpQe/Cr5gj+crkbA3uz7csRwXgGFPhC
6/JpvfueJxhP61u4hvRLFw9MN0QyKbSg++tye3d5Md8BzZwCFKgTvYAo0+Ecm+FQ
hhhfTy6HgVR2ldzOSOuCB1jxQuoHCSHRyNXwzg2wT1ERZnj4fTwUiLGd0vc7jm0d
h9V0gNmO/+ziJKvnHrz7lIM1h5hiUuAjb5DjOenDFsgL8kpN+80QvEVIV/gTRs3m
3lXJu3w9jd6nfv2pWC/xgPzDRBMlu0t6wD1SQxRDfiBNfWXRZYrD34Eoq2rSH5sK
2LGjksdWnvythwF/UbxnO+ujDeM1ocwPcYjaJ7qU4ivA98nslElFsx3qCzZSV1Tx
sjfz45RkHeZxM4H5lL+wCzu1KbA7jZea/U2zSZoR+ziy9rzmMTwrrUyN/den73iu
ny8IRkXF25xDJaRr8bBm50rhVJ7K60oOXDkhF/E2T+I8HDfSYoVCELmjVCsjQl5i
Q01SClw8H1+rCZPvw+AGpn+8rc1+C5ja5zVimx0LbCrHkqomTQPiIU94ZPdBf/zz
gwxVCVilDWetJZ0TnugAsM/4kMMzSVX+Y+ioUVchWnBbUUJRNebvo3oVgB/ljVAV
UmQtjGDzgY6+wFBNfyGpZcEqcA1k34Q1Mw+UK46hScJ+tPIXeOcWxBLOE6kKuQ/8
gsyHUte11eDGRJC02ucLGboVglzOYYi5QAEawpI/Hx+hXkaTqiyy0hcdjpLI8D3C
+4+uZ9LQd6hhmUkoy41RBuOCRC2S2n7CCXK8SxB+XvM5Qr8l1AMpEyu24yjAOKSF
JZMNcZ9tA0IX16fo2OMhPhBW66y2JAJsOc8NFpq27f5KWkIy16aBO3U//Uk6b7b/
wfMloLUf6uu58vonWFsKmiGVeYSdK0CuxSaGlzgwu6lLskNEoLn7Eva8+gCdVeJj
pEa85Bc9SkiZU0ZpNs3FmhtpALUQMZ6PkkZLZlAW/52YfBmcMckx/0zKYWGAD58x
yLuLSGMI98SnVwrZdWMsifDYY97KBeCW0ClGwNoJHtTHMNcLv+zIIYdfe/n/JWdH
sHR1DWPzdPwuTaqLL0D2OwZyJVPXwSJq4tFHMyUjxErAtaib8uN1jpeAkXs2mb9Q
GQhFzK5pejVT2xwWpfs9EMXU7jgHMtieDO4dyC1AiAhx2ZIuX212PJar+pCnycNC
BUoJyhH6H3xM8xA/TQa5FsnJDASnBjVir2dU4O4kP/ukdvpUZ5JZgXcCSz8G+B1P
mnIb69pZgftpMdGICo5csjykUereL66S749zqznLJv16ItmOgVjyMa9ZbDPfpdng
TLfURSdIx0SnlCX2zEJTTQGDGJFhGcLi0063bV2AtfLXOZ+YLprfUvs22FogqL+K
w5uKp1EnjjkFfRnOnFATjSzIM7YD4cw4Rn3qtWFcmOYBv6C/aVkL6eVwrpqdvnxa
RjVwCFrLKV9ftVbPbMkTVECJ0Uz1CyKKh8d+9laR19vF9jICWW3bEqi084wR4dZy
x6U+8f3rrp0WYRIzQldhMPKxZydumckEUZy8I0vakiaL9z0Y9evjZLYb7dzL2kQe
NW8T8bMIjuZJeT16hgGC2XUxVCN6ZYyVsi43Rtl7eI0ZMeY5bx2oTptePcBHF45M
d+ZexBWH8APkdFDcY/9gQlbkSlhhH5HEQIjD9XgubWDmRliTHKgwNtpnOx+JRitW
Ytjk6WmkvayZHt0ykucs4PmWVTbu+Zb3CKMjW7MsXrhEWKvFT31ObcQW2S33xdqG
KkLcYVmWMsb10uQ1hVTA6+s/YvnTAu1l1ThUTCdGH/Bmo4fk3jGwHtPz+AVFW3uh
TFkZMy1645+AM1V4vMhNYxX08jkxjpTAVBXWq44chyoodGcdQzNr0Fzktoda4vxU
XnxVnelhQ/RVnzUElsbtuaPHX9C+MZ6XuVfGahBRIH5FkDjrG2mrkUQN8QTgACA4
4N4YIQnrRhWRJlg2gV4vix7Be8SuNKANunTgtibZtSV92TxzW5e6yqQzS0ejc0PA
TwZGIjB34vVR9EpBrBn9lgDPvIsFH5U9otaufJkk5C5LVYuoT/bBLHFJERI0soF2
768j1AWYFan3g4nFbSV0yNLuyZZGBy53GqwuuYXi2JMddby54Fqd/1vkGKQyL1bK
D2yjrRdHs1vqafK41bP96slEeTy4sqUO/InvlEPpMN1WM0NfHrCy2p5hByii1+i2
Gbeve6qRbhNfqUO4LwQvefDYFNe6ZpakPUA8oee/r02bEvPUyEsfmmb+L6entiK4
dKSBt5LIraEwtexfSlunoSdGqxrmvNoosWPGAhx6euEJa9i8legv/BTy5+jMhGpc
kgLNoUa3B6Tr5le66IdRF/Qjp3M88QiK+jRO5dHMpXPAgz72U/DUuhz2XeabswrK
UXzX+au909o1A1ZRf9kUxNZ3ij1HnA9uI9zmLo1AgZlzF+bGqCo0iUwCju2t+eVW
cyeVlzyWX2+k8U5ytdB8qi6scDw0QjFkm8PH14oo+Mllb8MqB2jaxPGDZjl2QYvy
3l7GyclDrA5hU8dlOgVYFVcaeAzRRhCOd6XnYwSANgKspG+Q3HQZe1/YA4awOR18
Jz01H8jHlDL2MxNUgH9dDTCaGGEXwRhzB7L4kc2R20iV77KN3fnI8CdztfLZNkhl
sbpOWQSbFE0cBDizn7jaC84qQGRboINmOvqs2NMMUkNMHCFSmVN7yfNvFIOhG5j6
NDbEaUSv4AT5wHFnHAUmSbpUD0ifB9ezrZsOKkywEGuDr2l8/FkPAnMi0649YYMd
DESr6svQC6q2YLl6EiMFLZF51+u/d3v3tVQ8XSoDbvl9t9EFo9oBYcazHxlVtYjB
YuQaexDyrWz4N0KJW0lh5N1bu+MP+ldt+5xl8dxopznKw+afMDs4tXYu5MPbG9pL
igPgbHFzepaA38NW6AvDAIsSrlph9Wg2h0sQq1Hmv5+pdybHNg/y1sEuhTAjywnn
8aulhbMJwEj44pEl6xxc7qI+EmWRulZMoEepGsRYRAnXrSoK9hdczf860lBIbBQf
4sLhpdqQtxOZFsDLysYPvXW4ZBgHtoE8cdvtgWoJFz7JWK5MvGUxVaN2WewXiDhL
xMyGUK80NQZUFiwE48vsyVbg+WIIDoXdB9Vu6daC5KLJQkGQJDr+C95Jx7MV7bTJ
1XyzzNHvPkt5dXQpTJTTDmra21L8387SsSLKN4g9EYV6MUpAcbY/oMblODQwD02U
75XC2MJt/rtAE6M7JLGTHo26HPiscueNXrZkXpLR/7wY1baHCkc9XeSk7DZR+xqz
qsJIEAB6E02gLwVdtVrYnKE77fKT9Fus2rqKpINheKDHwhLWjVbfgafVbWImLGw6
zmatfB5UltzbAv5ZGFD2krFVYKI7OQPOTl/ldI+/UOY2Tk8F23Tim5FaIXKAXxN1
GmW7GHhm/mEj3q5g8/RtwbvUiJTNItgecxllI1j1/aX8KAorPe+mbh8wv0f7TBqg
n4wbobw8A21FpEv88S7kFC7UGIs5SymtGeffEhqtZh7SCDzF5/kJOVI3J8p+MvmL
S7bEdhYPTkkwH9K8KyqHk0c2rLjDprh6++eeVV6oe5VUB5VLE80pw3Lh5Hf1uxRu
e3qcEPENFVPUOuPBCnkEsBNFeoBqWI12eI2HSWNRaXyy05eiZOgHzSRLDVc2QyEE
y4K/hC1vfQ5uPOPaKp89CRgW5hPcvyINc9i77/qNjPHM9jFL0Xv+shOypD3I5H0t
e4q1I+tFrG5ZvO4KNfUooxQSHvWCbdBg64KkXyGROuEVkTXpehbzkcwo89+/A/iB
9tPhkKoichm45XpRstmGxtWqiB892TjWTuk5YGwj045lWtsAK4bo0geFNsX6/yNE
bdphwzcokr0dQOLfoTQtL1D2lAOYUvbii7rjnHfsPUu9SToCKF2/3HiOgXBSdBM1
sEGMYaywBv2cZ9cYOmh5izWN2whDaRqlzXnUwtByP/mC5omlxzJMKhbkEzZ3UVhh
YDNxo0ZW5ItwtVPbM/db0xNtlXX/gfeBg3k5mduVL+9QZ5ogNW6Xh0yc9fTALjsk
fk8we3hqrioIktjikkQrrwkrOjVFmvS9T/CQi5K6vhjn8ZOlf7rPdLPD/TLbztas
SNDDUauzNXc5hy3+7c//PeBQK5vLQAHCrWKIZqW/vdCsaPAoWJdLYyU7IlPGsloe
0/yHq1AIiqbSfVz8jJQ8EIDtKWtc8cKimx6FgdEH00yDX02vGOTCgONlfG/a0vbF
hHmd79vxOAEQqg6BXJ6BHK4A8WOzbm4RvDsw8LmBEDRnzLvV9ZIxxUuWJlqGl92i
15rLBf8vjIBNAVkNoQRYw37sVcXWtjcQ21FhWyFEqOEh0G87/YSsZYl+YU4aK2l2
rp8Xfs6VIrFZOOKQ+GMTXIHdq2IONYguMAfP4SdTmVx+nHYkh5JReJtM3TnpKx++
lHfJxgGCOKaLQt4qwwm2Bo2vTRGYt8lds3RAFp/oCXgWuPfgMu76f0sc9kfuyFkS
9CqpGJlf/P5lywCox+atr+nTG5ltC0yKOF/DamLesimjxYqHiu2ZY4pUL8HcKQJW
zhs67P9SeJKzxGUZYvGoUCC9GPZWpFWOazVyfh2pDS7zZ6SAQXfXScfQIbIiVWki
WsNxrm+zMyYdbuhNS+ahCUAiorLceXUB9NV5chrl7gMnkB26TJGPwXaoC90jL0TZ
BEggnQpTaHgSm2dGQLnL6kIydwSnovO/AKKTPiUkhRwlc5WBmNea0Kymr27pwJbm
IKlPzTgxb6Lp6z3o6nlqu4U3g55/FruqPeRSJoi2TNOQsMdNlCL8gMT9PVinxCPr
F1G/aYAMc1Hu58D5uEydYZXeNSG7HreVTmYBgnEBIGyN+BZGvL8nJoL57j03Bx7N
zUfdR6H0UZtX4qiGWC47G1lRc66JKtYSlRCn1PtXEli7eOC6D5fwCgW12dC4yQvu
qSwdLKiAcKVUoviok/Vfh+X2lQ7clgh9jZ8oVoBV5t9/4FrCSvJ3Vz8ibODwh+IM
6pVf4qtCCu+QZAO+NcuwjuqcbVE+f3Hx8FJ+n9V4Q5dZTaHfHDgML/jbhGWlr9ho
gC6kPjoOdGQE9IixQIGyUjVHffWASgcy3fxkzRr/jYNJpfSSFD8aQH7B0qqSEX/1
k/+4xm/pKTRbNeGSIfMSbyAQlMbDHXIdYQfcoCm497x1HWN+u15b49ReR2R68O02
BIOtIdmi8oIYn/G9xEqnJudPFk5mbMlmKeSIRIJcDPstuxgcU87ScyH+tBvB1qiL
biVNigPeKiVtjxDwLZUnfKey0h36w2YRS+Ap6B3BCZNjyEcgqL14yLdAKxLWkG5E
7Rp6s7i/Xuft+0VjEiajhZC4dVFDc1Fg78SY7cMYzT7yJnlVwLrb6Z+EHQA3N1vU
zjdlRaFtFPbsLYvO4Y0JieCQiWj7e+weo0cBi+I+/vOrfiBFjxn2FNH5YbjBaSOx
wAlRPgGdDiqVRStc1Qt0VhjM3sRgJzDc/g7/CDvCFaXXxgqw7PBLGlwfbYocp6/J
vZqDOzviSdXgm8D8YXlY5eEcywiIK+G8OuwwNwV2UroZ/l8xQoxpjAwtHCTlVUyD
FvV9FWBtc58pbCA4wfmYtyoPkDt7prDelusBge+hjruirmgohuSwfddLSn8mkkAM
2LwyXfv3c9dFYH/vNv/ZxmuRE2505n7aQNyuc0c+fBhI3zXveEHE7nAZIWXqjiH3
WlEcrOcgRH7l382JWYOb5VAAm9HCyMUV7KodX7X0N2fgq+MTkqjNyHhdj4F+Ljzq
WtpsdDg7+Mx4yAJBgn7hYLH+LCwiqsyH77HhOVr14x32SB4qo2XnQWRnR3v4wRNn
A6N+ixDevOiFsgDsrTezaJqIpmazcOfeXu/FDIPVkx/FYOLZ+G9g9TnCh+GZ49C2
aLZs28QtAqFzk/KKj+thdSTr1w4Qy4rE/8tsr+FWpcrGO0VqctZzOv7Fw8YAsQ73
Iu9ufieD2VuPYkQJ95POKAp/heOUEL9t3kxKi/2dFtgF2agRp1xQ7Td5R2iphiyr
cqT096e+9wDuTGn/Q0dLWyPqa8UH+w4rveTLADc503q4USuSE0AYA002CsbNltmt
AYeRUAbLUVSu1T4mBTtP7bWFwD09HTruFtmK+kN95Ju/XlB78uX6EO6ZnBnLuG8P
h+SSoL2YNrU7KPwyzS8zE1g3+Y5+wfrRQLvju1+tpXpY6G6t0R8iBpnuMAItlmQZ
cCMT/txQkyAbq9Ci4Asq6yTK9mi35UMGmvlvbBMz3cdXNTBmKbYQPhzeNKtZrHzV
Atsbh48rWDV/0wJNB1cTgUVJGySXtCgE2O7a0OA8I/wo5PdccBo6z7wCHt0zCck6
Wd5JH4Z8BkDHN9qzdCxHCcHMge/7eyEij70znf0/VG3LIQc+nlkxEaF52GzHGYZY
DIq+oUYH672YZ/lYKwHQc1OP6+WTldn8dtUxFTKtwSGJJSKhA+Fu+Kx5XTeMqAcQ
dHEyCcnzuZKp1vgexb4G3Lzo1SD70nGKjgxpYSOsDY9Ivf1NjU/sEYzFPx1+PtQa
AqWAxsbE7d0oIMmQpeiCzv2cilfKQLUdI0eeuPrTAaivEhO4xSLt8FUYrDfGiHxa
kWhIlp6UL30nSzsiMkUDbZWijja6ktteWakYTvp9OEooqsOucEDNPJq786bl/SGg
QPXjb6B5kHsUpWDM44olqw8lzjRsEfTKxXmvddOor1eKBE5z8nxvrazWKQXpcLx/
8noQQCh34Tb/pYz95vZghJKW1FdjzZc+YeFv1U06hC+bvt5Tb+BHyQ2ERjFWmqvT
qZ4aE06JNsl15jX+Az2YF9HmVsCSZnfh5rYUh1lS/pr16IsN4GeN8a3sMnvNDqvN
/5F5nFdo/mkX8Cxa6LbWF32aTEaSBGqYNd9pBKsPWXRu+YwODSCCcrLSVkZPnQOs
JeVDNGao0BnRkQr9Lxi1tXFZogiJUcuQ8003PfGUjbi7qD8E7hMQit57Bn1ywqI6
tnXc+ERPLVGkQ6M6nEoHZJ8G840md/gZuxV+bkvhqfiNQutWg8DDIS3Bl+8g0gkv
bnQN5KiCIWYANUGPy9GNMdnuTZWpBWgBSKUKo9BBscv2QCmlKg2cQgNIPTjjG2u4
17WfBTcWgAXGN1WkEHZlrZ5lc8rVFzmuTdck3ojhWimmCLnGwQOB+pRte/Yv4TE5
F8mE/WR5urJBCYy0C/cfT4wlNfauB4SLaxpM3uHdqi9kyk1oWhOBrrlzhfB58kBX
0zn2BZgaM909ljdFYS2zPFjXwJdM2Af3AsqbSj9RzJ/u3GOKFfIof4exuM9PH6Lk
lq/Rk/0sT0FHTEvinXSDeIGDuHUyu/QIZhKHVWoS1JsPuvC/qDSFE/FMB039J/o0
nvLjdLNc92Lvwj5pYvWCcMRaUvDQhSeRqDfG7w+vI+IDTCc6XlXj1XVfl2EgQ6Yx
QT9cATqqIF6Q5Xwh7JtrGj3zU9IaYqaRQyTuxAGUs3iXSBYX+2cx8OMZpL/TaVZV
fZwozGFt9gnulvSMfB0GuTVJnIwtvEunZJhI95tIZSo5Ku2GW8LoS6fu+BNdkUMU
JMux1BHQtMTuARE7DitQX4sUm6a36iJKZ/wSGc6wAfsFdBRoNrcv/8BhzcD/HMj2
zAChk3pfytvHkTrZdmgO/piiDgNZL7DghfCyl0SqzNElI28aN7DjCkC+Ri5DuP2T
lDj5cxTypchmGpyzEP1P/CF6rNjdEx2vrs1Su9rYXvZOBctqql/EIHOsHJpBWA5p
D+lQ6/ScKEGTfK1xn3i0KH2ixhj22+y6OYKZbWIaI8W6sYaGxiDd8HlNA8jYcVsv
IPXqY3b5/GusFUK0mLucHZIFscnXVajOloXaNdfcp5y91KjddF31n0GNGBW79krY
ktKc7RCpij5ZM3spG31GLZub7nzhWnprwZkOJkRsdoBHO8IdIpx1Sd24h0t1BOJV
hyHFy/uzGaEc7CeQNjCLOpJAcHMwLNehUXbs461KHQZ4arQ6F7Ug0t5W1uPZsrH9
ITA/Vqhw1J5r+nEADdJ+WHcB5tAaKiUmyxR2XrPISx1ylfEuw7S+Y4hX+ZIvjHMY
kDCBd44E5FCkxXQsSAelBMbXEOX3ArMUS0FR2N0OpWwHcI/ydM+ekkGf/GG6tipO
TfakTFDTm0w16hhWCZzizE4wO7JI9kVLcdWIZiZag1kgfHjPyigG9kOcWPImPQUe
5/Dyt9JNA37uMYWfc7VXdJz6XqDjPGdq6oJhwnAYlpJlPa1SmuzCBT8goxGDWubL
FypSLZ99niwCvsDDUXisqXPKr8LULnLkxI+WuQ7ufKvAcMvMeD56s0sRGPbo1slR
/zRl+grqTm1N4btoTotSVZTGkRX+vN040OL1ohgIgVy0lPl+douM/yn4NjOjdO1H
QwNm7CAOd8B+bgKOKet9II1SxlwU0UTjaJRQxvT7/2GmT+Aed+05Hdy+RirPb9Vy
kLVFeXiNEfbqwn10DAQgzFUNUIwhM8r34WCxISxj2kklvP9JDBUR9P+8b4UoUeqf
fDpwBej1k8plkCIik7Iz2AFeCAGqtkpREYxXhV8NSXH2i2yVCNGZI8c5nfJ231l7
azt5WDUqZ6ecyevLRSNzQ7v7VK931bQTSI3+Yd0IHByxswSbz3bpccmR/ms7GkYU
idO5GYnyB2Gyk8bSBkgzp7sUe4GO5D7WLlocXiJvG13QHRkAz6D6bC8WK4kbQKUg
erxTTYD5TvorzfJPZu17ScgRb71a0iULE/pccM20NIQTcNF0iBhsSq6xA9vXRIeZ
64Y0W8ZZEare8o91fikPfz5oDIUH5NWnQGrnZTcZOKzo9Ms7/7dcURenpNQeSQWo
ly8sFzUgeeqsjjpIkm1eMLg6hA0G4tWjEx1AjgYM8e9Uy6/k+5SAgS9pHyOuZm2A
HVudGnq14Jw7DszjNTUxUrUfo41w83oxkbOTVXQ3Iqh9BNalk5sJRgIB783vpwOQ
6ah0McSts73W0TAXXOH8ANg3Z2bLmz6NtsLeBpIakhuSxo2IfRj8xsx9lGNFoTIf
9UjI6n3HfLDJvuhWjcFvvBe6ApHbgxKM/ePIi5sMISusiz7w6Q2mKeREm6iXEQml
eUvlxoQJsQzUn7SeERxzxCG9syCDPAL256yR0FaGmbAFu7Byc4HikVPkjunyU7SW
ctpzpS7k7Zf9JFVMn4ly7d30ziQAArcWuYbaXN1xoNIEmWtqvvH0gR4f5twcw38Z
o/iI9S6tDf3hlBYr0HHhB7j9GcgGIaE7F67xgoiBHNhRv/Rq6p4/HwzE5YOmcBdz
rqtRzqJNc2XEaCYWKGYr+fDty3JYqJM6wCSsbaYsivKVkB2bgvE8jm/qrnN2ys8I
UWm2U1aXjNyeQ5BpQ9EYlsy7NBfxjj2Qy3aJJi25aovxdmxnSoqkvP8YHVikdleq
hNnC6rrX+LDe1+PjXgtIEnzy/riUTWsd/gSCAUbF+mb4MV8l3Z87JpT3l2H8AiQl
T97XJchVl9lMZTguftQnkwmi+x2VFcpRad21P/s74DqHk2ymKy926Kd1mXCtw/tu
dlnx9iv3DUMGTenMUnGhDKAs7cBYWJomNvEe78DGt+KMJfu6vftUve0MjMZLGC0t
frjbWva5xW+gkEKr0kH6xZ9HU9Vyn2qdSUfuyMkGbT25TIxA68xbLbpdNhrTtrs1
9lfDCcBYtUQM2+KOoQuRpQ/qwlvOBxm9Qkl1ogrCxoNfHjum0LEt+m5J7Nmryq0F
ZfbRnF8O2hsBhyYcOh0wE7AphfiUUlhZJIBIoo+d1QUwUlGtIaBs3dqjoB8C76Ea
IYSMa57l18gLfKMh7R1D78y0lR07Oaw2BMXs5PW+WUYorWuQuJ6seoy3IoLgUvf1
va2eBbE7+NtvuE3gsUEjH4OASCejWxxGUrsC7mtL22u5/swg7WpIJjgzKimOvb/5
ZekAysi8nYr7bruwAYuhcGm3p4cwyFb+LmIxOGpGdZ+TQkpfDXATJyKO2T7Kqu9i
Sw+GUiMBkeFZdE2g19/lsZXgVC+l+siWxZwM3gYIl+2yIkbT7C/WNXfLuoAiCG80
Uvtz7SIk/Z/0V0gt/r41IEqW933thiWTXIjERK+whevHuwn2YmvDDLfzj/+cBOlE
vkbnvdC5w2nAsnu5VGa2PZdZLcNhisj9lr5q9Y+jWKEcv5NFZDHdXTcEpt6+uOSC
FS6xpb8/1sHGpIGNXKpoigxS2OgUoi1awb6+R/wWuDQXybRTz5XQTEJUxlPYltsM
b4QDESvNOCgPrRftLk7ayg0DnCWD30lmbOskr9TqHIMVkfAB8rMK97sEqbwcD8sx
UL2jruR+whxXIR9BfwhwERuniHnUF5K0Sy5BFD1mrLRXP3+VK67pn0iPLuwFSCaX
Aic1Smy8ce5wcgc0d6mhYWb7+viQgbHgLpcI6uEvSNWig44nsST425sZusOoMLGx
E55wtGm3PJ3RmOqw4crb71CTKR89E6LIDZzADjbn4Xov9HqmdKgTpdDYmaY7HYFY
oWqsma8qhr7naBlf6EDgeH0YTbhgmgQijNp0VqD2JHtKMR2RWGk/FTWVXj78UJLF
gj6Tk0Et+V7w5oBqR/eP2VrC2JrQrEr+oIsK/IdrERGWGNhI9LLuqpETiHWtWuYk
zQ8t994QfP/vqka1duBvNe38VzEcvI84cPj84sUp6k974jP6+glCJU/He+5726AU
ultDYaArvAOYLm7hkO6tukDZJyXvtVTudY2BF6C8Xkam9LoEQREnCKwVM5dMMk+t
tY5n1CbQ9Y9G8LpmA09Id5/GQEHB4nM7HJtjXVkFKTrdCLsZOS5JArg9LM66s8Vo
lxKSCSmzbaHJxQH+pFapi4BPDBr6OyEf4zs80yepo3qWFsWNuljtCEkP1j3dWn69
mPoWBaqhc9D30TP+w6NK9ZazvcOilrhiX8+ljb0YUaufhwE9VKvikXwaATOMRYgO
gUAWjksC9CAqZgiV97uXqBcVSYC1avI/Ydc8dUSueuPxsy9cRWhL/ddS+lzP/hr7
limNWpC9CP3DIlSIDVjy4EYGvWPHFFDrZ2g6BOPQjzxUkc2OTA2qxUuMO7m/r/WC
FNCMSm0ei0soZKH/mvTJToWzvRYarPupZ0sgqVa2z9j/OsUPWdMOUmjzF8yUDZOi
x/+kDW48EROLygG9BhYRRjhIiWq9qB2lP8mCh6zZpVs9eQLalNKiebD1QMq/a5p9
XtkGjv37+6TiYFtnQIW7Ui4d+z8/HMpE93NseqzII5VjfGn4PWM5Gm/ZYOF+Qpzv
3NYYS5sgPKOoFw2zgYAGVgTmn62meOsie5R6PGZr/lWlpLJ6D+99LUKbUY6rasp4
r0DQ1Au3BAspIb7AGTAu1Y0AWvoyRSIHilSMpyJfDWVoBehhHh3JVPmDBhzE+hD0
DDTPlxEyftoT7yznc5jECtY4Jr+DCymHHXKYKAj2LJVZkP8wV6qhlCBwdV/M7EbC
yamH65HHnUKQ2FiildksgJRfg5rmd0B3al3mqDPiwHRIjJf/iWM1eo7l8MmD4hgb
1wv7xuhrZJRdIRJebQWHt+i4Jr7N4WOMv1mbs+Y+VD/UbPJUj/8blKoyFfv0z9Is
pY3TrOkfWVFVSXjGQf4tdpmPF9t1ntBtSSIVvKrsCPsUuBtDAlJqEHbcXWzNtA6T
GbraJhCkImPvyk+i32NezcrMbQxPaxebRqGrDgNiib33hkAIuMIz3H+YctAx+lSd
VAseFt9Jab/yVpBA2S6T4NUecj78qKnux94Z9Fd3H49UTHpm2BuKqPQFXUDpkOwJ
+/CpdkrtB5WareJPXp/jYmHfUFaHSlxnQ2Y4d3SkuZbhdaYnCoaDdlFLgqjHGfLa
Jlggyas6WWKrbuPwMr5g1uGv0mp3J6rFxvO046kT1P77xKaIK6fW2U7DjFtGSX+X
uFMZtF9bb9P4txsARveoIwECRZFbMQu7DiGGYstC8vNb8Ddo6FHF0oxnadSiYcwg
ugz2RlN00yYJF5EoMORuvcpwA7VeClM7tLimURcat6S0X9ro2bK+vLGfP0xtEW0y
tMDCvk7dM3SwmF+VqnZSfhWO2m/8b6RUkETgol2i5+ec8eaE+3pk6+bx9RJrkHs6
tVndjT2Icu4Z9D2dmMeU07Kvpm6bCa245bbl+F7iPMTvfQ7SlbuzEJCA5hmbKDdC
hjvi88quw7Xlu28XqzB3CaPhMmCGUVRPNIANkBwUPxOV5d159CGfO4F6b2QtAmzU
5ZXLWdYRddV2kM48yI1yx9Fdx1hTV9M1fSqOSxIL/uyJqAVc2sY7rPL40lxYq1pA
4IPv17KO5IMmRcSpIyJK1VtYs6Ca3+USlqalDuWAa49+aO4H5Lmi/c3tmUPn1gDB
klPkrt/qyYtdKy8/yr8nK5raZ5XoJBTRq5x51qQdPkJV6tlR3oU0ssY5uSVqzhOg
z/+NkC2HQUp4WUJor4n2fy566p6yGrKOI4xT2KIKkkOpNBMPz0nMcNau19tFN7Z+
JQfHMynuEh3Mml9qktOlsm4NgXwPP+kvLPtzBwo1Vj5/vWM/IvhZBQQzXyCh8zds
Ja9uyexhMXcUJVazVWOtPKT2GfRI+mV8XTR5LqaZUGuGlbRWcBKArk/9ws96xHpF
yusSYgQJ+WEKuoSyQyUubN31gTfTLVZrST4y+WXYsAVopr1QueO210mhe5jDoJGm
MLKpqchNeV9fTC2tUrBF/uOlXkWw8QRSpCN2BB5baFRDACJlJ5UDV+b2+3SmUEx2
vALWo8sk1QrHUm1oposo5fqR8uCfWqtquH1F590mPaN4XtApnCujP+qE/fgiOblD
DJFSacB6htb0mJ9bEZua5MAUgWTgLV3NoekJlZHAkbHRxRz1SXbyKUmftH4qSPx0
/cf0F6yDHuPxI1x/HRHMa+4YpnPd8Dq84TmKCoUtRWM9WkZDqzdGnKcCCBmfds3w
Yw/0BbwM7WWs3tzOaZkR60yKcclar0OZPbmI38GBGSRoGl+NqzKjnO6bQb28X9Y/
r4v3QJlmps1KFwDwS5zv9Rq6amYyYwVAn5u2iOGl7/LxPegg2VHGEnkjUgrP4sjg
K+1n2DgYvXochMQHjuwfDzzbZGxLuvyLDWQVIPpHH8O/2s3YuuptWTvyqJlCuAuO
GZijVUezio8vyLPhEGG2o6+XiqF45VKmKjACxw45kh/W+1BHnMga1TXobWnI8S7n
ZaGLVYflxtTul5/s/yzo/1xKwiJ3FmBYV0oP3jQ+k6DEGBk4HLcDlWjWz7oYSdNb
nma883YcVYzpI00pocclf3JtZv77S+TmhIgL6pO+x7Wy7f/RFYqTy2ky8/qCIP8O
uTfhLnBLdAOfvO2kTFyFaSiuRYh+p5US2uAe/SvAYyhnSAVDtADSzEtr1s6sfqIt
zI2alWIaVPj4tyN0/L0/XZTCUzRYVLfkgLoQhnvoXB/iJPXRFKH+u+gRYqocCTuB
gJEyJP1uHpMo2NvGxmpqA8gOYzwFr7ojXzFyqZwns0wltV5xX8BCYbXN4BtzhL+N
BRx6e3TX0qGBPtJyK6oocYSWFYzfEzDtb8+BIs4iGRVGcUI/ffiKqENFjPwpaph8
+SdANaWXdiHh31NIQ7s6YlRVmlOC2oRVYKfTVlybo2BKJS6X9zvXGDTpcvf7RAcn
Gzcqwd0HGYKX4zbzKlZqkLvgVm4P0lBZxBrlUihzogugZYWQh8LQoVegrHxXz7dY
Lp7rnifw5G6UENLkNJi0rze4X3G9SgHiAN3DxlCTBP47bPV0IVKWJ5Lh85LZs0EC
4tOIJ2oAl6BngdUAuPIdwoZQuHrnCWT3JxVp9GmPvJlyc3qVYEcpTePyLi16duVT
k5ugFOEatQUCbaJ8sZKsTMIsTHHTSJx6ECZcC5/kIxDkOuLeU0+FTgVfLgJu/Avl
zHPaw9E2R/rMD2rQcWFzMzEtiwYRnXRsFuJsP9ZNnRHa1ijDVVBI1XWC8ln7aQ3n
L5AGEP+4dljrdKRhsa73RjrBryWMVT/mgNBZxe+DaxJqtTh44qYXNzOqlc9SOpID
6TdPc+wP5QzFY+uDgHLqfu9xcMZQCREqiD9PW2WGqU0Mt6KEY+62XLjSifA59W/9
jdabsrfUakYr4a3mSciLx9zDw/lHQ2FTu24jhOX0HLWesF8YvfkYNGev0PdYbOkT
yVZR5BMt1fiIkD7qJjDV38GgP70yXHI8CLarCo8ejQbthsq8SOhyq0yGCiUg3SK4
Y8TDB4JTwTVlrBKGk4nr7bG09OU0xt/Z3mYVRRW+po0Po0aJ4wgc8ogaEvEALh+h
yUh8u+90HZ4owgRTOLf7JPUnP+iMmwpzWQ8HxuVkCEntwLPGUjrIZIe1k5KpJk+A
oLIGyrgyKkQllSBRcz6hxeulOLnPyIgMN0bKy7Pkd30TZe6c+e1/vWhHHB66eT7E
XKfhd/McV6K0z73bd3/ayyUpBGB+oZAmeU5c6fLJ9XufKGt4fTnhEZkI9ZATzkGK
LJGQV12KZXyBqIbgl6bgVrmCYKQaNecx3p9g5rSOQDQqu2zJ90GkiyI4FS0m3hlu
dk9IE6Vj7eL4nKv/It1tVf2eRKbM9dMeDfIfA1j9ZQ8IOUgT15hdGirPvkvTIilq
rgDyzLPtDhpAgzw71jfe+GheFJn8IxWvqtkEDVd4LEm7YUn9bUMkmF6B0FFGkSX7
kqohx0qxISH2sZ9tlb3GJ3b+bE//VQK8FO1/EJ7Sga//sHKatNKYxcW+QusLKZfA
NB6mPLkp7baXzsHbaTpv0GAYQnIHXW3mn1x7uh1G36sUr+r5+W8JMPOSQRZG+gza
1LkIqI/HAa8vJpZPrFtNAX5L0umtz3JDy8q0KxL4X5xVuwT2x5qzQ7WQNKgXv3LF
cXixpTdAo5s9XE0t8XmcZsqtBibHlygj8rRaSy1BFSSvPxGy475m2ZphCueuVLqW
YB1q/Y94V1CvvT1sGf3AJ/RcdYmvdkxISLduosvOCPoS7aDmJR5q5nzzhEDWkSqy
uFxn955AarrRuVc9m8GQbjO9ZFLX8oo8r87qwfhhwm60pNoPryIx0azkQwhDDPAK
tbrw+Bj1ukZDvSwc5sNWNaB6ipr8bCKgu8ImJfit6jUSdYtnnGzIrkKXy+I2oih5
+m+l1YTzBV9bgx7sozKBraK3aAaFuGuoTsUpGnEB0oa68/yjNWNnfN56seianFPC
QG6lffOs7qd9IvX9XzeE/05CphnZNEgjCIt9oEY2WRRDGM5Rx49IwNjf5cjeu0WS
vbzlqABEnSSCEPYQb05OpvDK94AU6bvfn56lFwbN4X9V5inz1zBLWm8kLWLlCEaM
vsJG84sxCNElX1MdRYESWynskLyDe+c5gp+a+3DFmoFIfcUCFlywZtbKAefTiSOY
7qhSh2FYNGV8L5gs2B0cdqLXMRvsAsgtlWl4u8IOhYnpRTNbaW4jJQkjs0P9rtOU
mgkFkvixJ3wfsbEF/yiX0NU41StYuy6+EG0EixVBHR7+1zS4QqNNqY3oLMALOtJZ
0gj+xKzVuGXKyIW/jisxzNkUYHq32RGr/+ETBdlbbtv0YoUtVcLzn1ANukDmgkHP
D5NKwIWAQkLoOxjqNZsDkmU7C7aKGHoqzGUUYp/bKBfh965pNDOt84hSqnkMlq1N
os5kdv+vlgOtLw2DjDMwQzhqYBL+lD4ZOlP3W5JWjVICdpLv7dX+AcQSMN3BOCKu
xJKWJ8bfl6zU4WDXZ4j4GhWhkTmhBKunXrrpYS5vzGYJYq4XN7sIYGCaQMddcmx5
4fbF1XUbsB8UccnDc/21TYgmejYcq3Ks0hv5AgXqJX2vNa7OICVtdgXob3rISfJB
zfZNZiDPHgEbbrmzMOwbSExCcpQPnYxCyoRXEX0CtG6EHqWen+J9zREnuXWoAl13
1Q/sRQn9S3R/uAnpkFoM2kDBPasVtwCrKOVb7idB35rhRELlKfpD7Iv935vJgkCK
AJlaku8QcUfj3lb9wFqs/K6HGWEQg5IfJXaA0m4GlCa1SbGXG8qp7KbWnOF10tkI
Uytbs0+l/Z8M7OVvZHH2dYY2zIVl2aaG4WRE/0QrUdKQq+dl38ovd73lkBkiJi0x
1pIDVWlNqyWkuuW4TUZYgplrlS/Le14G87e7KofHy0qysZy4puqtN6fIMmV2Dd7o
h7N7gLTrhZyvs+GtcB4LdV5k2VXMFQ4KiLKP4ol9RS8RfoXllTg4FCc7g2Pnq/lk
V/OPBgoBjJEVH18kTzfdGzJxohESNRnv1/VdfvsV385vEAGF4DRgIW5770/lmU29
h/ihAkS+OR1qmPa4BfdqoI8ctwpn5EEmQ4TUZkVp5LA3h8FTMJ6op+adROcBv/sj
nO1GTgvP+hevHtC0z0Z+bIp7kr7gn7q9Yv1F5ymkP/0LkKBUDJPinyPQWFVZa9HN
8yL1Bs6jvEr5M5euttPa1OEeQ7HRQHwQ3AJ3R2N2V3zq261NtzI+1o+09fuFI6Bw
wyUynqWkdNkFvhhsvrTYqL5ro8VqDuNuPdFjnIoxCTKGhCB+/laLL6aY2N71zzc4
TUSS7g2xKbd1Z4MmbDyzyUpGa0CS6bd6Nm81CsJnZxUuMGxtcWnx3D+2FLdJ6uk7
fsUJGr4ALB1Irqbl5VVYFaI5YGEjyNqd8l6oq6mxC1oMH0ghaxZl+sABtCMhkll8
l86sY1YaNVzy5SfDmVWb+kSgKid8FD5cJM63O3zw5IEx+kO6Dv43/n/JSZI0N3JI
i5XvYSdyWxL5bOHefFYX7z6m80Bl+LmQDV9D6Wo13BLBhkVoBby8bNmjg2KrE4TF
sCTyl8u+yF+R+HdL1B6MRN8dt0SME9JBuLAZBA+7EfBTwOZgy/P7P/wDiSddUJIU
2ZRv3bRzwGyvb7sVRhIVIV8qexSSgtkW2jNjuJHlNW/QEdh5vYt3We3ZRrbnhpxj
X/NDW/CGHR75BPhidO5GVUGQKVs52AExFyIVtDcaxV8WvvaosncbH1bHZY2VIhfl
iogqJwEV1U4wl6Ys8TJZy4+kYifcukJrc1+u6ypgf82FvDr4RICk24IRghOyPO99
GBY7t7ih+Yio3Bh/q1vdDwUcDu742mbylLwcoxqf7zMXDfP+W/Ke7RUoeOESevN+
AA48rg30pfcU19G8HqiDtR6qAmwy8XrSDPxx85XTJWVvZU8Xgg8dOgS6GCkyf9gv
1WhB/2Yw+DlrfSgQ91Xmqpl2jIbKoWAKx7peS28wBdCQ/J45FLUgdIgXQ1hI3gpG
DXH48b9DmcHmhw1BQHl/BDVk97phoxYy8tdRM94GRZqOUZeBKl1fwyx0sAZd4ytn
WAUrNCxFwqVBBsLuDfM98QbzUygpjX8Lyajs5l731PJaiVkKUI71PD0m2JqcCnut
cSuQMtlrSPWCZQGGUSnE9eq5IvKGv0NJZadg0WkvZOA68wuqdQviEMofIJhwuDJM
TWVbPFk2nBbl8wnREaRKBxpANZQpfaxkRgQ7M8o2cnk6LBD2onixvkqDPqlLwxFz
fGlsoJfxrLkAssMCnsmE/b3NWK+e/lukjcfl/iiYROCrieZnuVzA3dmY6llFzcZJ
skO3320u5R+KFodNxcI4KNOsEv92ES38PNzpe8OMTGktEQQiGhMgPfXkXx/mveEX
HgOOcRLIeb1YyzxY9Y1AxA+gwKKwgbzaqyLSDrCrvIEBbpVRx9lk0PsKSU1o8Tc3
RjdD5ac5CncOx98jeMPQRUW4dqzDAvWBKFTS4AW1qc0uOCunhBwmPe8k7i7AVYA1
PPjREeOxF5OUQLFKJvuuKfM06LZL+327pCO9Uy1y3z1+iWdVTwztVKuA1okw5Ddl
xy3qq9X7nAHqWuPG4wWxxubHNRam9XJkChVU7UCjZ6DdKfl/ShmUxWz9LozhYrxE
IvNs3rVaSWbNLcZGRR9ChVOooZLtvSJmlu1vpB1E+IQWLa/9FMCw5cr5ptZxNLvg
3LHvnG4NdD3HkRn8HkZyAQqgFaGGhkLaqInN+KqtTKbz+3AXt70LYMNZQqoxek73
lKShnSN7XbewgX1+caY47fMukKQtazfUG6+Dz3lGG0gQ+tjm8YoLLz8wmnbAhKEc
yioUmO7y+ObIOv/e/7QJsR3yuSxOMEaxZrMAVZXcsCq5sJ6ebVoidEv8brl3CfTm
mmGi7jwVrC8SyUgRA9KZVRwDzna82nlgRA+CX0ayCzwkvUNDYiibtCMugWvTTwWF
wnooI0b6JyQ935aiVhPdgw7M+IJLqINpiVp83+xYXVeDX61BVmguzhjJJSgGRX5K
9uzQ93WiWwq5HROzb18bE9e637yoEuVr6RpGkZbUwnHsp43PN/DGxO6vplkE4ypx
rcsCeupTqmbzXfqomh5hrSE1hShB+CgpA5A34kvl51qADjR+47LBmNjE6Ew+Xr74
s0zwwUw4wc61BqE5MPDdamSgb69OmSSjPwFkX0AMfZYAl3Q0gTfzC3QTxADgTGc9
7tbaqGCYzMrD5bIjQIJ4h7ek8DTLHPawkzsOoYpNB7Yq/cYkGLsjyO0q+t2WRQL1
gGS5YgdDihEC+55dYmXadVucDHoVtxWg9IK97YGltxKtK1FG5WBqv2nrKlo2M9Cl
U6bH/55lpc2zB+4N+A0Jf9MBpFHF6bs0sJF3S3Rj709EkZ9fZpGaxr/H7hweT4Ih
NlDCmFm1gvFgS+hPOq22ZL+nCnO8Ihkm7OIMumQG0GeJM6eKRNf+GvOyPTk4QkIx
/5sj1rJ4bB+K4k/5PuXrUumi+kOfmyJGWP2HtdnI9HmOrqFaoewzRVm/JrYNPb+a
GILG4BUFsY7qs7svEpe5IJgrszRJEnpfzBUCdsJbXN8mLM172Nl951eKzcm3UCUK
Tj51ZpjBqFb1olVScUf9BIuUn8mD7WP6nmnOup60gR1AeoFKuD6j9rH4VZPAkd0/
X2DSHayHGTds9mUSHojgiWm0NljvunwB7MaPpo1oxG4uA5X/GIBIbyYto8AmKD1x
ENtT6ErZnCabASpSKAJjLhB4OSOV4sK/n6cjGFYrqiXeBY0A9VIbs1mKkEeicJX7
O8IVy59EataWr5YqJ6ASXgjyok6slNVigVyRcPzx0d5i7u1iKasSmTSaZq3QJC8c
upaazamD5epfWKfxsjRa2ZBei/M8pPxVmST7GDITB4CXbCVNx+xHw09MgXlTvQ2s
eiZYOLO+NwVURQvU3vZtGLj1dYUgxeA+WFhNxPpgp167rnrPE9MdH1tUfpFWEy6s
NwbRMBm0ftyk9T8YL/QDW8lQ9hDio9eR5kTIDHFWNQqkH805VY15tqglad7mHTD5
wQA8LrVAc52MHSXPRXFvbshYHLzUJvofEPaBHCfx6lOBtnmTmLBye80PNYVrpS9N
dROPhwQCY7u6utrv5Lb7yhTqh3RFm/xty9vaVBDa6hHO0PxsFrAMaNsXaec6C5sp
F9wf5uXp2iwWjAyxhJcXmK2iYg08yuGnHHbv+Dk9WoRYa/3Q/korlWDWdzNuCiT5
ItWyMjCFUKf7Feh8sAWf4Lsj1B3SgQB4QDzkNLFunGI1xUIJTvlnvs7JMvlAxKyO
Cith77TV+aBlVPNPoYds6Wh5StKHDY4KQmG5+kTLlgdqGG4hvOtuk6nUjT4kVCjz
72WzD3gXoNsRxjI/pNay1QzhsYzvGGJtqosmuv+UtVBtDxuxEZgoq77qmJD/v5eZ
yA/IoEJvtFpJElnHP3HQe3GfCWiigb+Ks+lME20QbJtHntY1kMn/mY7d4UiMcjwf
V29aXJCpkabITNNKxs4DRLEVe6qeQ8xGNDJ7o1nmsVr+1MAOp78lYaUHcgTNuJBr
uDesCsX4tyK/YOf3eg+xHnlEhxkkwb7uLmvZVqwhNtyJzZGktNactAXev3jsmSHE
Kdnf/aMsq5Wu2hNY3QZ1dBpdADXsWr1QS7mf8f91Nijr3opiOb139bLuOFXrpUTf
2jTLkwsEJqVcmmdFmYBZ2SXTTB85uha5f7f94zUcY1Y3Qi3jo7kWKMVaKa1Xa3aR
G+3HTvZD18JkvpxZEF4ViQ3cF3dmIOVZ0m35TTvLF9EgVcIgfdiKADaKZZBAjz73
OqxS/9KlS4wjsJ2HxhOO+HDuyiHbBm4DuBCDJko7EShSMcWrxNyqalaTz8ZfQLa/
dgriWUok1wudQNns8ewq6fT2O8lD3JKvA6gZyCjuPous31Dg5wNDtpc4oSKa/US/
XLMqc46mn3eUbppm6XfLxi4pSpBXJ7qS/hiiKU+hVPVMAiM0uRlyypaU2Ye0Js74
1D3xuMrRvy4cGmqCNDR4u4ck4dkL/S6oLI7vGJP/Bwu9aI2Z80ErFNUc9RgF1W3J
2b2hgXlStDTvC0tvA9Ls2WNu+RA7njb3LqKfZLpja+ylNEqwunUye4LV0urv6ZpA
fKZKIofmI2MrRLtkmHEiHeGkRHfY62/waVn4r+qX/wLDJ4bDkkwjqnCyqOOJ41q5
qwRC3sshdfD1/96/nzTbzttrwU6yVj/0JUUxTeJtDZNHpNWtKqRZTOWMp+SuDdnw
e3MLwftwrbygBPIq1HNhIa8HNlFO1CRbpu3A9Q8NT/VrpZnnGC/3kbTjgRWH23e/
QQ1DxBqC2umW72oCldNdsDWyZ65CpyWR9rIx5r/1lZq8C/1xIOKLXTwTQnAnQ5d+
HDMCZ0WWNv6HLBx/a4nfYMIq2u7OdaRSgXoamPU6iqJVrmFXM/r/olZQSsGDgOPX
RxBvL41UvOwt78Ag5D3vNJsApx2SoPN8mTX3+gl33aq8KxrucoBE1kXCRwemiWzk
Vt29zya1x6a2z82tlqwkV8XQ1TTBBikeGi7v3TDHltnTKNEmlaZnGPNpXWiRNXma
8w3Z128mgCLjyK/fYYEu+w7TGEatabNgD84lNf6oxOKGjpAOoMA3Y5hjkS+OsQaI
Mk8B425GTEoJP+UPFxgHPSV33wprb0309emHoSPLi9I8PTkes93hQraol1xt5lv/
SlEJUqDSiCjVQmyefRLKrCk9t9RpwceLwNVnWtyPHUVDr0usoapNbJZ+8pwlyqmN
Ms/p/KAgEZetUo+pCSsy3yfpssY6+OjWBzzV5DPkw/uQLHArxTxV0hO+e0TmRwMM
q8h130RyHGcchqArNA+/EG4iGGVzHERnOqPc7ke2nz/YDaOjnt0Wm20RDZ2v7gpf
5d3Ef1e5yl6iXKNVMswp8hTFyr3V0Iecw9f79vIZqs9RrNvOliKFoaj7Dob49m89
TtVRjPw/UEXLwjauW5G6salNPhlUwDY8d5E6MhXrICc/imkVzynlj3j3i0c7qT7V
b5fA8RG98+ezhq8i5w0r0nZdb7pMEPSq8TRkUOezYl/ZmyuEfUd3uiD4K1ElkmFB
6VqJtP+uQgMjvKld/sFIAPwmQ38MJdd9cpIs1O3sIm1+JQoAPiyrKWSgk/n7E4Ka
OasSCPYKuK+5+6V3GYQNhkny/j0X09BM+chH5Z0d9luGYAGxYYxSFv1YkW+xb6xD
wffXGP7hD05XidlfnRkdeuqJcPpAaPqw1KGTbOCnxTQPFf2/j7elnGKZ9zFklgUB
zTy/KSD/I54Y3KKNY4PoshpSR3crieE/NluYvOpBenook/AMb3Pdwfg73FEwGuPV
RO2E0pCnlPcOOQLXhkk7ShrS1h1OWoLrzXkLwkER+yReTA77TdST8TEOxcEiP/RP
BJSQj/7bA6awqEsMJ8kjzE7BwOW2upiaEAF0kVLS/VZ0SSTKzi0bCrBwDb4DOJBX
NhBt83maMcs4qTH1BAVhLI9PFl1AkQhiKhOKsLdfPYhSzAzSqEs7LkfI/TcdwWoT
evIHs63S0o+wW9LrfVpGKpdy8qjrHu9zp7av+Em/8xX6PkDrJCk2WNUiVbenCLMr
Io13ylbDiQhv75V368jXc6YIbqy49cEfixDZ1S5phaTDCP/sdfhuZ1yJ1bhInE0F
KiZ6zpHe5OUVG9DZzPb4KE+Wfjea67o2kDWz7XneFCEQEDwXSO0sXgNNFi9eF58C
rQaozeXdGep6457A0qcG1XmBUq0lfFQZCJogzQ25feEMvhu65f/mdHaYWjqTuz7b
bkN2RX7r4kf27bdyjFu6YFOBTpZ4EfnmFaAIpgrcRv8CKnuKwAB7cuFvXCdUTHnv
VD19F5SYcfMuS9cUHkvAguRoESUSU1ssZuwafAcb28ucHwxcHMNJjfMAz6AXvrr0
Hq34xheKsFgjlHC4GyypVrGOD+fNp0HCMN5tmyTXd6Gi8Q9nEjvkFKL5VHBB1GgZ
YVWwn5URN7hiQnUwyu+b6VwOgO/o92vWyT7ubGAh1Xp7k3NcJ9kw5APeK9pHJDZb
6Fa3XG8nQNjyyf7MsDNCYvrmHZZkPqv4N3+KXQyK/u5Q5OX16Ufn6XVKtB3jr65R
1GYyG4sPIrDP7KqAMojfJ4U/MBInMkDdB541EK7eE8fdJ9opeaU/UKgu4q6RNIdP
Vj4eydIGm/HaadVOz86bILmHyDIjO26of38mlV451ea0xfTKVQAns5hbfroeBuJZ
vqfqbiFTRQHdOLH7Uv1N+sautjfInv9Kf72xV2auISwtpisc8ibvJxT/ZcmzF4cx
4LUjoKOkJlXAUYB/faokRP1Hk8eov0LnOzGBSlVmcvgNQHIQ5bChjYKVMXDt9Nxm
oWQ373fVa6JOl+aCfTSGl5HdVhddp13euhgpuX5ImVgFQ8GdmnStDSJWcoXU6wSv
eYdoNdkve2NEk18W32Ppv0sP8Mez2yZLXfxW6stDA+NxzTdsmqt2P5qSrp6Pyxro
Pr2NCSCOYg7pGWCSrt3un6jvrgMxXm5ZS7ZyiRaLvHdcW1eqYk9R5bWLi1ilu6Ng
MqYJGfnctAwjOQFNG/603o6TtlQ/uhxq0GL7cGuvaxqMRrxFMa9fjiY/z8d3pCOL
EsDAnNVI0hsJ/pWo5UPzLiJ9jKyRk1rGDfMfydvrI9qatRUwL+dm53EmEU++oKI8
k9853VKT7fF9xLZp+gUClvFh9zSJ6Qo7y8HEb04Pdr4pmgGk0B49P0oXMdQI1nhO
r/c5S5yfFr6FKiZxeuVlEq8/h4DFr2uCUwCjEoe7SE5KvmSstfuMGeOMbaX1Pj4f
jBi9NdvDHrTMYY454kjmBBFOZ5kfZqXt1ok1510JQ9P6FNrbQiCuQL8+IfHRU3xl
B5++AFqlwGndygLGGxiRNZZ5KJmjsAkfRCvkK+H+QSdUn5jIrT+N2wV4Inesitru
5UQc3y/VdY1kSo5jMElCzT6Bsha/hTM679XOt2BDMfRZ4RJEC9S0J9PCawyDZvfU
5paWeD97SPZcaFbDijjm6ddVJnBpdPeAhyOZC65Lq6ey6KcSe45aE2E8O9MkpA4E
XMSOb3n+xtcdPPlgAHOHBolrDTw1jKmNfOYQ4JOZk16bPayx1yVrSW8bX1RmZXVT
JFUD0CCysctCLDpqORCPlbhkf6SZhC78sv2gqdA/fanJFWKGNbAO/Hc1+T7sIYy+
rylgc6Voi/DW6c4xrufI6rIsDx5THQ+uT9JchIyJqMyTvr9aERvnLCOW0vLWtM0S
g8qS0Q319vNoaHi6c00wmz3RHQviguL0nnpPvQdBXu3fyn6jo/M4RV1xxUgAMXTs
6gQkUF1PqROkVI2kysbtwjaFAuk6xhs6h6/wIM704wql4jglppkqaDslmZ3c141L
ERM9L5e6PirAQDG0zq5UGpQ+K4XFwfWGyCUGB4CjZsH4y3HBH02F/fMOFbCC8ag6
cMwffe6EDO/3T1ddX6CCVWfAe98Q6X8IPivoC70ImPrYpiCA+jKjZBsq7+Cp7Kv7
HKYhfw0vJfyH/1Q3UuIWYbkEIc+gJ7PueFV2CD/7lZdeApCvp/XAXyYrszz2lIuU
yoB77uRgEZQ16kz5ORruVYQgRsi8TcP/sMcTYUVcqUOKWbF/5BdytM7VC2wemo4z
D8VYFS552APvJNJ6c/MxkZuP5OHIrmZqL+UusVzzhcbSss4hPJ/sMVRr7IGU5bDd
Ntj0Ypi795/4FhsDk1ySvWaKFo7AAChsO0NKQVt7IW8E5IjI2FPDDV6F46cpoLtW
TvGrzeM6yvGWmihA3wMMuIt0nkG26FvNsiu8PVtmKeWpDGeuKdj6JLKBAwE7hlP5
CpjtHdcW2GZptKLyy+ji+Y8hSxwQ5Obb8St2NM0IKOrSJjOM+9kEfDyc/6yRBlqg
axO/3TtPT2uKVeezxlNr8PV+tE4GGXqv2VlmLTkFOOGGdgkDmOAx+LO8ASMEM1jv
UZKCIdHhq4tFebuEsusWdeZMqg8+z2qISES3BZelTx2L44xNSceSYX9yyFeTS6nk
E2nuHwlkIdqy/YUt/v0LlVsv0x0vFh0D/z2YGes9sbGe4NWdQ2CvN9NhbO9hyCjU
aHdqEHj3/y+zoVdDDuBxeuONkeI7WYHdJQf/XgxmVIzQ+SDEjCdTff6q3QE2f1m8
ZMEk1z0YR6BH58Na/Ct6ZBegYqvqR/tGaKPqQ0RhFTAnlk+LHzKzhEYBvvR5PayH
F+WKS8quaFcsBKFYC+/QUjDiveFncdpR1X2ghDtMxaU9guQyCflIL/2UrQ5Hq+Et
wTrabRrMyP9SvK65NBgrUfng944XQfn+nAY4o7DlrDUGo031Shi6F3sDkr1vYcQB
l2KYDF8XEVjkBOoIqq1DVqR8iGttU32qXc/yc+KVrAXE9h9w+8W/wFN5pF9ESzos
og/m41m6lLILMc1u69qHQVXFOTUe0pa7LrEInikQCft61rC1X2LMJZcGiEe9zLhT
+FNNUVj0UWKhZodK4N1LxVXG0EurVTTZ6FohvISdk/VbSRJRJ8m1Z8NkAlwUyhyj
LzgENegt1nxVltVxPRYeyBGZaAXzZXiKcgjRPDoaFnI6L8up4MUlBqlxiJKcm0rV
wLRNwuXeDhlnxbOq467uvuXNNQj7ejAoem3JX1RcKQcZIRspnoYKyluqaJRRfQM0
xrJDWee/VklapvbtRLeUm8rVEC3VmBj5M/uyW0tH8J+uSIP/LGQM3F867S2Hwm+V
PQOJBKQ7fV3MGmSE6gck8tuB9p4+Nmjq+D4E4rKOnHMewqlPqUXIKCo9evi/iCap
3aeNv6reHtnx6dPLv53j2BHQmySpapBqWB2ZLr+/TJVVp38Rf0v/jxWJAyTc8k/d
gqBaoBvRQSbgno/jKLKHmP8ULWYs+vS9cS8HzHUoZjUlRhjUdEuEeQsOKhgr5us4
qNmJD34YpkuEPnC3RUNytjz73Spgmfytlpe5LJv12lnhWb/VKLP9xc5SSMdJvU+Q
t2nH609TCUx2/49uqkUKE6/Axsb/fxhZ0+Vz1JjBgEzpM+jugC/6j3xzNbz0dWjy
Gr+BR0hk69k341+TlmnQCDn4ut8qWIhC/95SIPI0ES8jNYqo7Y6YAeIqY4QgaOPn
TF8kOdcUjfqFU9BFKuXHWCU5qbxm5Zwa6CyE83YrtvCYTHFlX1sAXaMlJfCfH1hQ
e96p3D8Zi176DchhDQ8BzDleLLdJWSoNNBUE5foGuW5S1bTpFXgfghJXPL1Jv1qR
WyuBfpMDm5oGTmJ5IWFNcMEQYUgQ0pm7d+aZdmoweK7f56kOJgjMOlJDts4r2zTk
NrK7daz+QaTbwEn/RkfLj0UNzUVCE9bJMEpyq/RxlSg0XyzqiPV39VmakINSjQoo
BHPMfo8tljRjc/KVNJGQJIOO32pwqzHugNgejOp1q7ydgMdAXez78k4NM8Al+CqE
wJI0bwT1g7MLBcEnDlnvIxlZ/6SSjMcH2sgrssPie7CKsDxXyhOWKZSLaweStJRo
0yNaldvl0oqD2DmnnIdLSU86VUAxmL5S0R++Th7jpZMa7GlkIn8hNe/lzk+vdIyk
QYjb24reRk2QDbXK4kLD95tVsfkrAjYBpogDQuS3uu4cCvGK69aUrXSWXX8XWpLV
2H5nEFoUnc8NZZJbJ9jGnKLdVcHG+ba3rSep+5C7NFPtEUon4d57b0boAZy9SV59
JrvA3hbRxrBH2HurVCqjaf/Afa3TudDc/O1/EQ19cMsPf4K7TMbbeA2vSn1Hg1Gw
TSxtuCwvOSzLRoG8DhQMVAL2XWMBR7IpOjGOukMpUVe7pBEVzYD2/Uvdrqa7E/cj
/ZxM7Oy8pXaMHZe/oBm7rRdzV4OMPx3MZwRU57WbYSE7rs2SfG/NHeowtxbo6vmX
zgkbQpXCbqJ21v3e2Twd9rFWS4H3UNA5k1FwDKRDIpcs0+nsOahi9zsCiJRKpB17
cJgVJpmEzayrbMVocG/25iBcP8HOc5XVss9NUR4Ge3RrUfKithF8n6m5zC8vcU6I
XBrXkRbsmOY6jUHsA8kkeLIiEqX+KskkyrjfMTC+4LxRpWCMo8YE02KBdESuwyj1
hBPAtEYlJQnZn6KuwTEeI4Vw7VET+hyci2L9jCNs6J8Y6O27RgwS0Jpx0fifIpHv
PQR1wfwTGzO8D8qFcyFRXfGYc9F2bJtfhliUc/49KyCUGQjplK/DMnnZhjYVLw7w
/1KlVZ5gvyqsER9+c+9S8vNwDglQE8yNh1akKZXtqoVU91dFA7A+//Ripjm94ke2
/XpRjWMfm4w4LzWQTI3r4Dsc/QdxJt1nz7M4/cNi5DdawWk94CXW/6JIlNW7a8W/
LHc4xitMxMDaW5UYoC72jWnP4hdaGhim+rd9ilRTSN40ILA8cnlIV99JuXUo0Ujy
OtxcJIvQHQuCHq75fwFQ81GYLAlmHmZc6Yy1Zvgg6hryfCkg5ErhTg8TIU1x8C1z
JfXn33Za9cPpswXbocJMewk779mVmcqgTT4Ml9G74InxZOaCZ567cqC8/vfFacGZ
8Bh5SVCv2vOWqOJD9yT4FsRGO/qLWkjkIeS2HrqdbZLcEi0OaMC+0q+aiUo/0VCT
96tXgVO/GBADPakEcof9cSITFRRHpXPSbmxkHSy0oQ3Qlh/Y1EICZku0WXtdIRgV
GjiduomXTpc7+pyt9faIPYsK0KbBfCPQpotWjsvBX97swOxY4q9CiQpbnK4fOdE7
RfsFNakbtVY0mkDx8sZLW4ktDhBv1nbOqCBPi27hr0kZ96fwz+mN3T4Hv/HfAcYD
jWEvNgQ3/Xm8b7fwcSRX+cMhEDbPxieMEAAz9lLaa5fp0LwlJYoJDUQvThfTBqam
pVYSyN2PONRYVqQ2pJNK3BeSGY8GRnZeovT3WqlCBTODysdX8ZKaKh75yqLMCdop
q3UWUJ6bgpSCu1mtDc8cYP4Brjj9zAv+sZvMVnhjjvuY5ffRKZWsIXYP1dQ+pYit
Z1bhmABUFdK+qBmZOYtpte7KQ2PHzRCXNlDzakeEN6+Wael4QmwvUl+4MdldfBXv
LOzv0BlIjsOc5o6v3mx+HfSDT25MULZbQSGZKoZqS1XAsUc2eQJ9+SxKRlNX7saS
xzLFIxHRGASvagTzVzvRHhz1tYOKLf55n1a2bC9uQGy0YYmLCKQ3cXbzKSnjOGh7
OKJzZx3JS1/rCGka9/ec2wZbL2tntl2BNjlNxscfCRrQHo2+boekpp/c4HylGo+W
t1LWwBbNyccSY1D4Ov57ETm6BWK0u4zTQ3ZTLsDuzgDI4PgtuSd3gZtN3xcczQ0X
PCfzytnM0XjAPch8bFcsiCmuQ6ui8odqgK0BFIz0JukFSxMwRl02pIq5gzaYfSHm
XMyx0/Tel1E/IK38BgLVy7+LsRqEIkbY/Ajinit2EaXMOAXS435RCHsjs4x2Yz7s
bVahSjkW9jAKrswYxhifIdLsFirDe3wL6bJqVPsFBs8uOfnT9FM6+C8b5BJ+AOUM
KZ6NHbEL4ESi0LkGc9PVrLh1zWML1yXuBZ/5HmgIi9TuuDQdegE2SsEkhFY9/h8Z
Wm/5+Hsrr3RBItpw0K5/4JQWi5xRBSY/rZB1WnoU0MsFbTZBmfZvd6g6Cb72MwV9
SzLwoS7sflfU2xagMjSuEVjLLNLo/kzSre1OHcLKYv2NtV+z/fgvupWD0TeVUEwN
jMvO9QT7q8LHH7Ko+yujpNkbDc8G+s0Jz9H2GUgJWGqB9dWThee49lwr7Hzoz6Ln
BFoSxH45vOSfESbOAlURY6s3SbNuA+YFQMJoJ/FAPYPCjwE0gi2QTuX+8xKTIZEz
Kf90IIezF+gbrBjv/f2WBDscsWJybNqE18H8El32vx7/HdCsK63yyJ/9/OWpRiyq
e6SE1+rihCv3sQTI2qxM9qf8JOLUfm1F6O80ItA5JqXXU+AQ4n2bwqnHCP1H14Ur
PhUfrC6mfcNy6i7SM/gg3OaDRiMx+VA39ToQLTxJfvU+lVYEX8R/YkthnCSNBmvr
sRyuJ0mQf3bQeXsAJOhNIjV9KG62qd4yR2fssNQcG2vSK+x1rhCyg7IFPWHyXR5Q
xZJ13/Hmttk+HygVAjCRwB/McHi6dfa9UaJxoQ6nfZXbGy5YlED9cjM74o3z9bxR
L6LVK67IFtDtGMnUrGoeIEye7EmXKVSVO1ZnmC04DnMawv6PmsduVdIFLfVBgLBn
WS7NDZZhHMBuuwRBQhUFjH0GamhEJTpCMdfBQIzC/bFXPEoyHmB9zV6kWpu4gXM/
Y2VIFBOGZYZvMOQfY9Aii/q+FmL+8h3Pd4xxkPf53g2bS0BKG9zc/AZINYgZF5XN
3uAK9WIEdAECqYZlw1ztEjAVpFfu/azIidYGBczmoNu71rDd61TwxF/12vBaVEwy
spXMIBHwtI4dTRRHRbpI6nZXfDMDvgAN+VWSqieDGYBlLwPoQopaBBiIQPiYVB8X
rSbLVRkWDHPWDTix+1PwQQ455lIIBrxQC4EEfundJd/cvC3ugsFN2qmVky4lznI+
FWy9iiKTjs7LNJ4mgVNrEvaZwzomSaJSuo3CBmzE5+/Gyx3zvN0+URjH6oAwsSP6
YzcQiKrGBScb2sXgfiB8cHwG8zccqpxoAfoFwUiVSOPTq7h7ZEBksrkcdrd4a1Nr
cZOhqBFxkJmEz65Cfs7hgfv6aw/hkjk5kIUey2YdK7TglL4hWzQ2YMFNefAZTBKK
9lPUddQdpcTZbhodrjsQ4Ue3+Ms2NftYoQW+g2hf9zRHFOc+QCK8VWRoYOJZv2N3
u5eUfsClbIV42+j/s9esu/zTYImQWl/hd/cRqYvqf9uy3362iJOqbrnVDJvoXVeD
owh19CItL+JKkWBGKAO++4t6mp3dsJNiBsz2naklgLDe8z0RMfFsA5HPKy+aWgEq
SpPSQihgPagRHqAvWW81bu/5lE8jCwh2zkzXLhlTf6NrhlwX+Lgl+Z6/fsv/mUA7
EncdzkIbanSWPbV0xiMkWIxTSVmj/f9edfAAgeRoMZb2Ts8mHMsAiE48AMIxMdMJ
RkpYESMMOk4Y7hRcjLCSQAJKFWaOZlCnUmWAWA9dfplNgK/FCVcQZSl3/fcostRQ
WjiJQN9W+CFJnUmB/FYdBJpEy4vW4r9pPb3+LszpxqEeZFMawYiRfzL+Hg8QBKUZ
rkYfaJ/1qVb3kgVrm3d2IDWthTpx6nujns3kCAdI01qkBpCgwQIWt9qi0r952b/M
5b3/e2pUNUsphQYZ7k/Tb2oTXl5/dYaLvgToatJQ+Mm+nf7PVtCRWtOdvuGzx6pw
owCLSi5Itnbrun3p6HFoYg86NROdAvmRP+g3bLUktZxYK450u1B7tmSJQ6IBUonv
NDTZ+k6P362pmTrB8EjnKAz56+J99hxzbleTI+go7drsKX53XaiLJrsoyEhuX5MM
uaIBWMGfPYj/e/AwGr4LavUIZsMZ9ZUaVgJw7Feydy+P+OcRSd7PeUD1oHlQ+cDN
BZg6R1O3HdxV+OWfNSS5UOYDA04dhr7Vfmm4t5Onr+Cq19//jwZJFS7nJns3oGdq
haW2aO+wHxSeqnDB6KkxlVPpVzxgON09BiyNySTJ0eQEWa/Q0mGgEBGS7F2+tUYk
ud77GLDxofffoH9rj+ZwPb211fSqhw2oTvFhehmcGsg3wMWvkiam7L6fVMminy72
EkXFF3nr2UcKUBnjx8yyX80wh3ur2ztOVhz/NYWN04UwVwO6dUMOa84u8TbqpxqR
FEvVT+qQyNbdxf6YhzJxA8SG3YE1JBQ0T0X6JWPIFzLwWVfzogeyrm7Bh3/e3Rid
OjVDNry7hz4IxUFsGyHY4F9EI+kW9/x60j5Yejl0SkHKXqH26AwHWrjPK7zvs6oH
71mYJ/DH+S6xYG11s7s25TwhNbfXjs8iIL0cv70gxhANetA2aUROXaxoaMDNXgwR
iBvQE9+FKorQPzhMn1lXkF0VXvbzrAhInow3LkrgWtkkk2LPKeBlbyA4M9IdPJ+f
XgM+7C40hDtxTX1NsZW9ZDzlE//xa+lLEVlYXDicObuQaGwB+Ey05RBoHIHxPLEL
MnOZoLvsQ80tVzTKcvbB9sVkK0+Ar4exq0qSILw7YdJsYcYPjMmQ61WHQsg2F/nM
Tnc7LW/JPgfYzVoTeYBQsmSlvoEW9jsXTpelbgStnVbPBwF8iZZuLdEfxY3NO0Mo
186GW6YFZTzSjopT7DuYjE0FoceWgDELDhH2I4/SL4MAn2IxIyCiNXd2a1pxj6Zr
HEWh0AQZc1RrkNkhWauzDjzHQP1XWAHIw4LnMU/pBYcaM3XKR+WFt05RU3nPNJYc
BeQdI8l5pB+8MKo57062mbxpEpH8jZhl6IWYAPrwB8E7MsMop1ZWcTE4PZLdMnGY
k3bJ3idU8FEK+27ZmItAshXR4kc0NV2AcosKvM6NLeW5YdsNtLaOR4XqqF9iY+jT
tX658fmEydHeXORlsNhqFEqTyKcBIjbR6xQIU13mtSLdjdkR6Uitss42JLX4xuFb
nFoDVLiXJ6QX4dLNKfcxwRGHoGaihQyQihGP30x5aE+xXCIMMN2PiydOxbdh/+R2
A4ZZJ2HFjN4LxNj0QEyYL8GCutznUrqdWKZezGaQf2/jRwfM1//axpQWsvDus/D9
2d4RZh18FFOOix5OIdZ3fiKaZUCoQEMwzaO13Szm6S7qAWC2VdNTjn21DM5qgHHJ
DYdJhb6a6DpkDlHiQh42J22Knd250Dv/vYB/a/Ezbv0jQeHqh4XnhMU4x24nT8A7
O3SUxFiQtmobzscG7bXWe1Q2AFWwSsA46OSDScy7WL+L/tpqDt1mCOJRQUPOLeGu
rtpRYZEWaF/A1pqmTI3wDwzEccUrM5pk0DBZBGF7v1dpXBKQzDLR/fsAf9u7jNF1
Z88+yXqpNKRFpasXa2H4HcEJwooGW82rFlFxf3krZ62qAEwZZokLM5e6ayHETEF4
xVgtQKDksQCZXns+GqTeIfn7BqQgYY13euvBFpM+7VCBLZZ40ZUV9oJZbwmmaXYi
zyx7roH48z08ufVYG8d0M05yi08snCDhlZTWY5JXVMGwAhL1nbTTJC3ViIUZ7Fhn
Iy5QMN2vHrljMZI4zx5t4e8rlJy28YmUnuQDjDwnMJ/hX5xMl3UYvxTkOQJZAylW
KEUHqF5U5MLK9rpjE9L4/KNd4NsWJNBUYctjjUmptBPkOn1PI9K5EV8KyhVFssel
nVLM0CYsiP/7m6moEPlAj5403XIF/hjTqkLeSLjfgN0fGybMXq7r2TKLlvhM57j9
Qpa5OfsHlItvJIdXQbmTk70peqCkS+AV6OYGkt43VD62dzMaVWShY+azJYRf/OLD
Fo2Q2ZgRfao+ZVDTzpT6BxRxELpuydGfVHmuNCCrKDQDrN5fRWyunHYHnfc+1A/+
j9lLi0ziaSFeQPDQieLQoE7z3qM6mn/0xABPwDWredUy8RgCqX0R/+aJAYUSJ+JP
DlIovodRSKMrsoKS57znN8AHUC6Np63RXKN+qxbVPQ/y0rOAzohWBgC1/dd4WyWO
wBL3ikNADnJfijQ88TcqEl6hySIqoL8lQRceL3+VVq/XbBu79CiwzQiJ1ahidcht
rnEWIqJWZ0A8L3r4Pp8s955v+4Wd+Upjug6BOzYnQgAxS5U3pT14hi9NuIZ93nIn
dAvXeZNP/W5zH3xKyE10WUrl/5OMg120Z7lM5m42EGDNzde+X2CT8GOEllcU0cha
fzLqZj+dncq9DCzHVmsZb/ZtYXUtjFrTSJ5utlynPT+RHrVawgVkcdinxlN97eHG
JiF48X7WGgbwhaACIv0TlAHUhwjeocSKWcfpbWqGuEwp1E5d1ASdwdx8KrDpoE6a
INC5CJWzXPtuuhmbU3SVa0btbc1TdfuEsLORgpIdLYTttDtvjDbW0UBa0TLXspH9
0FBFHqvvZGD45cu27ZK7oly0HD8fnYkfCvW/KMfbTVQ/Tr1++ehbVvwTuUJmHmkk
E8FzdD+jQrYqJAKOpPELYaoap2ms/JiMBbfRsotoNoQ2sZK+YdzIyHwowG914OU2
5z2s3wiQ0TKUpA3p0+DKDtLzb634hhSNL4kX989Q02hQJMM7J3n5F7ziQ5ZUF4XW
bW9YpL7Bfap8LBHLoHEv6mFgysQvb+L0R5M5uGUzMi888x0LVV0FcD4PbECm2j7j
CWx3fZlTJHhQjaWS1/hT/Odn2lbbU1DktiOtnxkYYfTNrBl2eLEieOQb2dHobixw
igwclib/pYFAXnSIay/wTZbTFLevPf5MmIzuHw52No+BbZ/5rqQ9v6fQM+rMkZJj
n9ADgZUZ3zVbTfyVheVM6W7kte6zZopDmDts3p/evzf8G+vqlm8I/lH241ejXFz+
Q+Coy/JQlcHHBvcv38H8Vl+27zgOqTjmmr0gj6xsYzNuqRQmSMCXh/FRIb6CWQKD
XqzNJsHgQQwKV+xC075sPxUiz7bi3VQf1ZhwEwH8jeYRaamlpsr9O2eh4cxnGFl1
ZzlLhQmfnpGeUW42hqFdWUBJo+P5AOzpbd/1EtedWGIE8+tuFjNfcwGg5vsQaibK
fcyuNgLMt/qR7emcOwqDMD4izwr5INShJJtSrvJ3jI6vsP4avi3uEIxx/HF5fW7Y
f6sbdbTBZib8dxOxJM5jg8FHFXF8/j7xlooGpsJAq2vLftVLOFUmkUYF1F0IgMTF
aOU0ognCg0Tprg069HcHaAK+X++zKkndPSsKSsG/ZTDI49ig/Tv3VQnvoA8PSyxs
gK9lhSCpPOD/ldCzt6Jz5PpLP6hcf9xDueggL2nfdwyJrFyWSVF8xferaaoOqL+2
elQQYOoUHNr1q4pPKnXdzX9QDhZsGYpmJeiTsumdxV2btFvMVpwEBfhn2snjdpfD
nZzSreAramGTptl1yUz3sszMdb4yvOq40+dhpMfCkDOyHHyTftj8KCzMSciCAGQG
CKMpyDXYAfTu292Pbke7y4hUbl6dR203+b2aWxo9CAAxVbiZHYbzzWi9lwURb64H
kppmAadiU1J7CwH/ATOH2jjhdO/Phw3zdljvtki+JuZ7MSkilInvhB3Vn4cirsrZ
b5wcS+hypMvXO7Md65GHxr+pQsQUPTOteuSY6mtVF8fXtVaPj0lok7hlNP8JlS5O
aS/uo3GvfwPMGr+3rMJReBAyKBPBxImpQezVbQ18lBgMz6DUQ99Kjuf51nE8ZfD+
k7KC720qA+9Le1G6xTG6hJ6WxKSZ8aEbRk8v/ug0T+9hHsR2kOyCsSB5umfkEPXe
0oZb0P6c/CkLIF5XbVnrYwtXriisXhjpovS+MmRW63/1mL4Btfmr+/VZv8N+xcly
LOJsc2li3a5S7+Hmj8kygdlRY+vM0hJNb8pFhmKgudwSr7sFu83KNaKOmnI5bPUO
RVsHuOapGkQ37ZRLfkS0APkt4pGlvuKntmMOzckDMJNVYxuh0WNihX7tXv1q+Gaj
6fLjlrGVC2VuXsuRt83KtTaeaGPArDH08FP/qD2DJUa1Mu+G2Oxso1BoOhGbziiU
1pK4LWvdqeJ85HbyNlCf+XfOpme7QHks0LABJ3kVFZcNz/iTBlZhW2k3wEXQ8WEV
O516nKIOGyiF/mliKTAsAKNnY3GhUsjjhd/JFvYtcVRZIskggJPb2BjP92XyhNoE
IMwXgVY4qSzrnKcYd2BK33o14k0KEFnD2F2YJj8iwQEhNCsC+OlRVgSQky2OiAwG
ODCVxGyVrPMjNQA3b/Ao7Aj5FwjTGZAcEwhAvms7cyOAxmVnW7M8cKDu3564vt3n
33pwIA2SrcKBKy7JbtcVEqraBweHn96EEa3LlBunJz2XOEfC/8yEtIIha0WM+/tx
Wix5dYALUO5ePBhWZy6z70mKyjNLyWddZct23fwm4zwESbQtSzsZ/zFBp9VQfvBr
cIb5aGQ1nw/M1MMJ6QEOVPVFeKi3cFIZoh9+Miktc/nIgXuUN82IFYY5jR6rpc5h
sZ+vPlSHOvo6avZY0LTC0i3Y4yP8A+Bi0H0up4nN7qYDuKkckkCIFg88/ogeNLtP
1Fp41TSxkURIcN5vPoZPpCZZCoaQ0KhFl6aZ4/HOzLZx52+KfkArr53QmupkhEzY
0sO0YyzHpVmMYSkzO/a0juxmVBJTjsxprBLU/ecxKok0asHuda+VUiXOAaoNrC1i
1lAx40IB/A/sE5zykq0dHg5QbfkM+SgI1XMp2OpwZhCFLjciXXY8gba4UTywstes
0miMYQDJp8LCrUD7k2tZIatE0VyINzt+j1hqMLIz+HfRTnIPP4Cj36UBjIwsb8XR
BM/G7Z/7E5tJk+SB49S2XM2Gy/pW6fKK601QgeQrWzTEBo88U0QwTxmzMcF3P03O
Q/BxT/aZlhStcNSW8kQDWGCTV92a9draS3UnxD7xjg3eAJ9lf4B+8wxFPGkK0j8d
nMi5QvG2U6tawN8jjcwb8vWWs+lfeO9NI5GqyBO4094hENKGjM+83+eX875Do3eB
6CNDtpv27Y0IdwWzvSA7Jh86FvxcgtcAr1/VhCxF+TaR+769GPSFbSBnyO3lq8eq
ogeYnN6TsKKMW/xRDqMqpS/soLf03p3KdD4XboFixLb2ZfoFcr7gA1X7tdBWw+Cy
OzdxkjEzLTd5g09N+FIaqpT4N1ckEUjVbfmKKu5IfP9baP437CUFatEHzKIT4zEi
WpUTkWb0zLsYTbj9jxOkE1qSGNwXc8xH2MQkR70eRoFRsLpIaovVeylQ/zcfHz5G
xpF8uVB8P1AYroCG1LubAhl95U2VdQihZ+6hic3f9Laja/k/Ex+frF0+X5qiMkN/
70B6t3GF/07vEJA2RasxwkYjgLeoJq9u+xyzEOh6t+1UACg9Meh3dBIHVXZkQ/mW
uHorWkCGUcTjRAMo0DIEOYxLCDlOfBWZtpG/ejoY9ze+72HphTnyuB9VvqfdyGR2
lIeUYCW/VZHtUEPSK7b+XcM405cowMA3e4/yM5ifhXasNW4HAQyoMxZPwVAGrip8
4UsLaiae10lEFgNtxYAKlO8c7NDoyeYg/yANRZrTBscU7la7obcrl8LDx4YaI3YD
Enw+e77/Lxf5GqDDLCWDqbk7M9UlTd4h1ohXevf0MA+5fSLClLt847/0J/qdMsc9
m1eAlLBB8pSuxtTY30ALwaTRlVDaE4R1ubpPYjdpgERoi7aaP27+rGqKeqWzCv7X
AvpFTYYjlufZzYQJKlH3FOsXgERLHOc6y5Lq+gNVAhRN1LhMi0PI9WkkmXU1HnnQ
ct5cgNPalbVTeb54X3O7dUB4kEPEdFZCyJTJJWONWf6uNPx2UypCpx5iFK8BLJ9D
xryIYvwwq6iSf6YkhaG4LdVpnNy0JRA9RfdSWo5yeSpyypLcbYmOIXdLr3jEgQsS
R1+85riPiPGcvCSmBKWT0eMVKfZKCsf5BiigU8uHieQWPApSWN9Td+u7Gb0oQVo1
0kiQtZwFIWl9oeirOAtoqRsHM19YjHesng6ZLV/rIebZBX6xIu6aUSrTB3+nghW5
wRHj3sF9G8aSmr0CHCLUqWrDbgfBOvTXCr9iBm/P0QO3l9wOHZsVZc7t0i3Rel8H
g9AD6tjGVkdPQe6RprOzISNFYgmPmKAKJJIJs0t2sq1C6w3ua7GM4wjYRtLAvf3T
SZn0SqUUdHQKCAsmehKXHbIUbTxdzupQGZw+/XmEJ50HYIXA7Okb1BY+6dKh2AnM
nsaCEK1TLGQ5jofr31KZIJI1FAx5smDQtHBf0MlqdXYKjb7dNsW+67pUfsPZ3vk4
rPFYFWqDK1QvBDaA0p42lSD52KkVGZzYX5XNdoDxA6p4sXQ7cUJYlc8M4xYtNMzM
egbYzN+sL08RMufBnPNib0XvrcbvewC/YatiTaY3aklxFOP9s3wResDYkMN0NLon
3MwxKcV8tf2fR1gt+YzMVmwuhxM1Vvx7CXzp0hByGacSEqsqH84uglyrFCEBCL2J
jQjppg2HP0FnJgRITGAO7gMQyLHXdEPlrbDzJjyoXYvUkC+bRzmtdUGQ7mVOh+k8
ptMK2NdOacb2a9HUIRDAf3SW3RFySBY0sVqZPiraGf1vT63zJOCJ5SL/zmnw46ul
1Ta8/kDozf0NfePE5Bpvbedvo8SluHvk8pWvH6WmMNENH5qsZVFgdFa83POEFTjQ
asyKwiaHdH1lUG63o5xyiCiuBkT3A+gH/aMWjsSRxrP7EQ82rOg0v+eNGdwNesr4
RkmPfBDyI/hvqEUW5u9waptUDimsvG8GKFh6Sz8+FFuhAi+DZrdtT09+QDaC2aRe
AJ114+SuegV+3YS9COuwveJW+x6sENHd2jcF75VTkwhIO7RSenKSwbBF1bK3Xqzp
GwsxDGoadMhQZGg0Z/ZN9qLtRbpfw3PPE8qe3Pv6vcbQDYefLmg1A985rdzSWJkT
LThsh8yNQ6ciuAskQJyxGarvFq8Q9E11eY76r5aqU1FstUfkY+mKY6J+2zlDpt8P
I/zqkpir0Ae2/ucpEdRi6CrvVINJh7Tkeb46GeTREEA+e3v3HC6JGvGhtAKjtW96
RSD1agxIwW9lRa4nO80crxmGhKE2BZDF8BS3RJhttNj1kj4NRhUmS02wgqR3gsH5
qyzl88R4Q4GP/QWysINRCA/N43+uvOkk49vnm1BqGw+2aPwT3PBEw5g/lxsle21x
NWSAZnGlPm+UKH9ZIcHDCiqw7G1Sf3rDBoIRxqIIp587V3pVnPaxWt53r28ZzFAl
3yFrbcbnQAXHKGcLM3SC77Kc1faYmgDqXgs6lCpsfM+PpCsyqwuy6YJbFRZTsQJr
jResI2GhwhpkA75QPI+m6951zgOulwHi0vcMwhDJ6VMebk5bplkYEiaEJX5ybTsB
It2QyB64W5eomNBXTb3gUcdC+2LzXrH+CE8J+rRny+4vkHHEMq9PsFDfuTxF+XVK
nFhG/PpLZ6IiZH+Ft+6FL6+C7O0B1YjKVyk4yM1CeavomFvxLZOJnk2114arknHb
WjN2BlgvTuHAkg6+NQ6jz9rLZ15TOhxg8sWwwj1FIY37HcABIz5sYeEmCN+lgXb8
7WOjk8a4aW0sXahKjz0eC2vYJjSioMlWxOJzT+fNH9+y5jheNbamrf7FHfT4ic1l
F47w/Ri6YzJAz3mb33Qg2nZdJj8p1fYQrVMQFqIaDROdZ63AMsdIfHmFodLElDgo
6t2AIdgG0J41pdBWmUtN8X/1R5AuqfGe8gitwmnNd3Tjx2J5RqL2tqAGf4vosP/i
Pd2DbnEix6EreOWiPUqUZS5C+He8fbab6iUDWFQDobnvidPsEJmuUuJRnk/Qq2Yv
TmkZdI3ceXz3w5VG5vBCS1lDqDsyugcqjzK/L6EcLDvi3vhe8my2rX7jiUrACevT
9s9ySBrV5AbJyBnEw33A535rJyOouG3n8LDwL9UItvaPL46xh25/f/KMLMH6ae1v
VTfjpJDGEZ7LRQxEhbBrIctVL4o5TrdcOtv/KY4TthcqdywaBet2r6urQEQ2iIjn
4hR/7ehg1s76gNQLadyV8S31YAZxwRCTqNTseSITnMsudPnu85LZgg/EQvIOLrvE
F7eqEHAI8KcuU8YEwhQia8ucJ90nz5sHzMtfPS4xOE3rzJVHlcXZKOx73eeoWq2t
/lebYu+JpvDR6yK2c3N17/QjmiFNB7XIBAPjDiv6+YHLQdxc2mcRQltSyoXdNQ2R
1gZuy1BH23LLiL+mx9Wm/G8e3DaonTlpGkgv2TC5MiNCE4zLYzPz9D/2V6tMsDYK
ltZ2G6GIC7dm9vhhRR0RaWp+8klEeJVQRCjlqk34cWViCZwgF+3mTayZTMc+IVZX
pepZtBRiEQopiF8ew5J+ZkbZmA4sKjVH0FendvHgyi7BA2TDtjoi0cZTzNQkT+Gu
r/ar/VUY5dWOReKKj2ZDPMZaJENadCa00OrhzMxrKnIrfgQc0e90a6m9aSjN179J
K9p+R4zZqockSqg/UmJazIVVB7ZqDzNDVGaIT8xAeq2KPjAcfZqedAdjhd7QNWej
UmLNGwZFK+Ek9xk3a4cDMZSul/7RYBARohHoZOoPqrgGvBIRGV8cN/7RQSkMLzoQ
bmdA1RqJox51U9ciMRAlJmkbE/OWMZxK96Kq6HHK+AjUd2KatdrCF5CDOIA05KMm
wF1SzYXOGbSRc0CfKkRweRZK/V2xg7/jF2oafOtr2cj9pF25FGzUE0Zh8os0BlUB
xXVvnW2/Qh60+PgXbsDBKKB5loKAUP7/RFEO72J419C6uveUTCcVZuL+CPC3wkgD
T8dZY0b5hwx5J33qPgim0d+iAvIvW9gGH0ivAAtijkoJU4NZhGw7PtoEhgVKBAUx
xjSD6EUsev52TEKSg2vsvFFDlkfy0KTTLLm4W5hK7/sA4ejuEqlWFQPOBUtif3fo
41nrAsfyZC2U2nBLwR7VgTYf+sWnGcB3gJ8R9CXpgQg5LBEaJEYVrv0eMKrbhju/
ZTMfeXbNiR7qLNPLPexDZuGQWdtwM4pZDU+OtzKWDFYnppQvJ/Z+v3HC/2JuRgGE
ZBAK3wTng5jwxUuIL5F4LWM3tdmxz26WaBVNe7f18kdTd9tQTYHIzaa0IQbHZ0EF
lzRqfSJ6Cv2JaVJTiiyO4bvrn8h0oWIR35B585gtdeIAHQG/02Sy9uKhYXxuuFm8
dj1Vw47urDFGJRFSs0P5OYuQdaYXCFzfTih0ZOvszsF05BD3M5MU91mgRT4arUbH
948I7sHYY7eZiVpWKWpveMFpRaRR8ivG41g3zCIM+Zybr6T2i5C0AzwlIES4bKA6
RIGQyZ3GnhycZ96IhGjl5fp4uzGxCH2o9GBvc18WwoLFNKrLpMDmCmBzPy1lTdP6
lP4RzN+gkV+RAwiKCDSSFm6R8V1g/kIDiCqdmREG1MicaK+85kTKasbJtXWxyN/H
QlvtEwQsJCrbDpz0YH1dbnU1EnohTrO+u3X0KS8hBuboCObxMdL9zzWGBYx5yPcZ
MZ5u97+pZxRRlTY6ffUm5tTHk4dsjwNNvcdgl/7Vj/Wqwlg13vna22GERTtkSDsQ
ALOsUBhslfwEvgXUIZITTK8IW3cSAdPdZMEz6+2Zw+CvocA4PkyA3420u+vURDfV
LvnMiZbG4up89RkvuNx+XrxZbIvxiTaC/IuiKdir/l28wjnwjuqlcZJPgcL2V8nZ
MjiqLiJxfRFV4xvsEj2/qE1DZW2U+1LmZyHwQto4D9550iLSoaqOpotS1rbencmn
WRxK256yfvlJMd+tMwgd7gFmyeByPqThS2VEaxhgUqaRjs++5dcBuBwLfO6XGHY3
aHK8KSqJSmAiiRHNhd0z2eFzzoFcqZrwzky5KmDbnKTG6RuiEojS3GcNqj3j3CDQ
3jHqtAbXNSZDOtV4iiUvzXP/3vJzs5fFpYfNZP77/FsoGUj57wVAjow+ts8MOXbZ
Apt9gUrba8xUlO5I95WoYPSXS81j2bQFt5wXanzzeJoBxMnFIWu4G7dddMBXlVPh
oO9JUt8oMAyRUzRCxq1AsPAQCLiLLxuIS1NCaNZVguPW39H3/qMx23uN+cOGm7fm
rbY4S/Zy1E9WFmPVqQztE7HAnFmOz10qbZOJ9aIOjKdJRPUSyHE/q9SiV/WwYkcl
7AybTSc96S4zrmNVC71RZIsJnxDPpkBkhkr/ax4k0/KL4G5i53ZOg8m7J3NGCeLH
KmDhNRZDeb7aybk8ccXqrr8rOxBAKGCvJHB/hOhW189nCZoIOoXyDYcz2MK5BBnV
OAaVgVq5+qdKvFEGFBQThOTcqWkX0zKnqXCI7rYGx2L/9gE/UlKWDTdtGGCTV5f9
kzzhL1vsK8HaV8+JVL1RikAjOoMToDCr22AH1wUZF7hOqrGemZco9PSdrHRxgyJ7
KiANuXIYemp+LUgiu0smyl49UMsda+itqv5aH+ukM4ixf8YojXiN4Nxg16/L2pFZ
NHZgLyh18CkIZdPceHbLLAMHk/RLbxZI0NDPMDL65tOwOBEqOAvJxOQ0jClxgsnc
OVP1Bf2qsGuMmoL7V41SRU4DF+ZqbrSC2QHVhQVjSeg8tpURKZsDjsa1vf2x64v6
sSVw3FVtTPxSwa/phR4vNpEk5/34HMX0y+OdqNVEr7mZN7rcvsTQqU6XNy2l4MJ7
eMgryzxzbQjt92GRHGqcUI9TNV74JejAE37lVRUg9nUjH5g1DNlkpLWXzHni7IGE
Y9d8JNw51YVe2mB5w6uQVcai193mCqJqyJX3BhNkVhpa8vSWhjNEsZ9SD+aK1+AK
e/XrGOawbSRHXlatp01leo2lDtiPflF0t/h3BAKWNaNJeMjuegdlF7Uf2uXJaxEd
Xji1RCWprd5T6gTfORyvc2St+OmHFxhsYk0b6DSu1GanCve46g5pCy/pwa2GEnyK
uTSl6uOzKGyFa5CBKLNt/YLrVoKUPvOLzfXL5/NS78q3z06++FE6OuBSOBtqYVVL
tF3ByzKiAmTmBmLAdPpd3EJfPbtAvpuNG3SZx0hKkKGC1r+cIwaVO0IXp4NhFvdO
eVWZIj93xVKD/FejErCMal157wYTactt2U3/NsG57QaESKUB06qpR/33T3MWAbPM
avmbgyp1XOUxJVC+aiR4HjTaC4Z9In7mmw5ZXdoo4rYaA6FSyK0Fe9G2tCe8D/So
7AOi1v+clzNJNFla617qBsc9lHzb6vxz2ZbJQWFv3lAJ1+mLzzruMAV448VJM1uo
OqbMGWQgv+XZkArPzns4mWayaLd2f7K27W+GNpKR+driQgxyaqD2qJu/Tp5dwauI
XQ9G2+frChRVS/AkwIC7bcKqxU08+Cl6r7WxHX6vWqzFfSOxPs0h5zIQJaXMmdhL
7L2o1kJo0Brn9yi2/Tge2nz9hbPCmbGtPAc7rPh5DuQFR51GkXYNLGSe/m528NI9
YoFhnKHTWF8PFX4zgXcAspUCT7KVz2eH1VSc1FzTFxlZ7IeMjeR/1r0uxxmK1tZH
X/EmbbcrKW2pXhBlr9VpcHbKTzXzxGjieM+vzSKybjP9NzlsSp0Hntol6jIASY6E
qiIV+LPA6YfCKgjy2xsejml2SGf/wNZB/PelHSSGCHsr/Ka2uyQ1/XxSfbeJGqs6
R4aVekSD1ts6wYXac7eX4Mmz3zQUszNdVdZIKNtHFrw17ElLIN3VXfj7gB154sBE
/A+ORceAYKQU5dCqZXjrvnO0rOOpvQmD6J5VS4JDZAGDtJlq4bCWNQRArjSqPO01
nDFIgH8cdFyX0iXr+KvOIExcG2GYV4TaEY4MRY6gQrPnyvHaZT/hx1iMb6pvTaDF
hvZ/vd64tJQlV6fDzC+5PM5ejnKzhxG9XPrZ1KJ8ui54k1Q9J4Olcc6ExOCE982B
JU1tdGEL9V5ERUUTw+BnYkHVMyHT0SZrQBXvH4k40h1LReNpaW2pqmgLLDsOE/iX
yz2EWrKfrGqHVrkQHV4FFh45nuGRvDV2sLlgRHZnXsUwiLIwwx8QZfn3A2J4gOy3
jrpXKubFLS2Zja6Bj8bekFzhc6X2wZDT1BG95RiK1a8x5jK5kVh94uvnOCFEXEaM
due3VycJI1gmiwZAhepMIsc+9qaCIoBkwUxkjB9GsZ8XFDWSW2MRvX7M6k4ICFK2
Te/QNwFQsIN1G2QW5M5ytFAeZwv6l8nmQIx5x23BGsUcySwpHh2/gIqeowh2fmot
sYdkbv8VDiyWPa+jFiErdTEVmrRGO/ZA0Aec2tL0c6JNU5nz5aw4Z2tTHJDvD3pl
nR7+hwm+pNIWS2biF4DrLzC5DxQTEIF2jzMwnnL2071bQxoT/rZxHDAyf0r7m5ep
qlhG6ajjlojfwCR6ZmPNK/3w4FT4WkeD4b1tFcZHjVuURO1NTIGNKppg85gEglae
1P9lTguveYhLhIjbeHGdqd0xdlzSFMMWv1O4ONbKJURdVRKw8pfm/Om+vxny5CPH
zCh0Nj7VyGh2dsy9993IC4zEvStegHkvbFz4upxhtDLO5v+EKnXCkwuRqI9jWuKe
Mhd6G2+QJIId5jMS8BKiZENwNaAwfbOp1yUnhu8R0jnZMsUGh03MDDR/FwnZDgU2
iucWDv0TDlDc9GE9QFoLhOoMXVBLSM/iSoLUQ3JDTGgLK0Xwxcn54VuTgpsvt86Z
pe9TxQwg01cNBuC4TyuvtSBFieTRJUm3p5Cgq0b/XCTzZ6mm1och1p40df9zUtSU
ffSQ6yUNAaJIwz3W/fzu74YlNYXVLWAovdbDYcAVKE68dWKS8kVdutMZTCKnTI4k
HaoiTv5ECWk3/EM9tJEMydcdBPyCW4TD/9bIEDpEbJhjlD3nGJIcThxm/NkMobRs
MijP/TA+gb0ruPdTsW15PtHE9K1KhTzk7IjH2aE2ohPrzqM54YP+74ij3ygKoQpB
eqVtjWyMJ+tYJpcr4LejO4T999PrL8sHAzJXzbVSUO7tzz6XMm2CV1ojJZs2pVKx
FvhtIN4GpGgRTdkGni7NnaTHhAiemuo7oK/h3uzD635ApOOZKfYuCr+Cn8gmrAX1
R1DtitFPj0ikNu9fN5LbWCkugcdP/lZNjpXI7a66WYfAe1hLiDPqmrEd2vs6+wli
vQ6S2OI68Mxvu/dsyXhzujM7HQiEMsxbk/EGihufrEq3Ipjh2qbkvMfqwgBAUX1+
ZmLOX77lxliuydGPyr6e+I+aA1t/owoPZnIaL25TQCTE2om4orKz0FvtOF3HqL5z
WpwWcmCEDo2nRw1PrdklWsHWxBZA8lYthu93rvYDt7R+5PtN1MWxKhQe4Me00evV
tVV9aneiM/Lqx9sNIKOptIAICMWNfRPFkBhj25eptGPGA5MshGV2ZSK7Hm2iK+UC
gG01LZqxa6fWqTNv0xs2hjbqOVsQogZfoJWgIQIxX0g4ge0pJk9WLm5OCJsy++2L
vpWlTjv/cotowgMLP123xzwaGkBmbTz1ElpyPdIpYkXq2eg8BAWBqoEbYGV7NxDw
/OyvN7ZZTV6WReMzn1rrsNdm0blnmrY9oIT0NensMJGHEKErDu/Qy4PP35A0Ymba
edU0GHZD0FRFXv7vJHtcBDrer1U4eTL1bIQHGerjb2LLfmwvl9NZ4neVjjIWd7au
uy1Cmyve/qEi8g3VFI2o0ILTEedoKPjk2+3sXk+6sp9bxBIxNLJBMSjkuKX4A5HN
iRGxUnzff/7KPqsUEuqyE1Zhw+5CfYimu6usvp4RVJHHqYrCplBz++/S+73S18zu
ckJkiFajvmXjK0s46/9Q3cyoMbnuHPmNHUVghZ3WVJbm8tAIIWKp41OIdxZPH5Gf
bKwLgD0BqzWna1aK6tyVwK8oZbBWogSm3Dy02lN0+kH2VFDkn2eY9Zjk0qdKJw9k
NSR78zlHEZjYaIdmOr1QPj4YKYimRkeHjULKV5OvZIE9l7VMSmcIOJK1qz8t2KWA
GTy8ePTwfPNI+mMO1JGnbYt8mJ5YRIVjeaYngOaDXFd2u7i5uaTqvoHZCuLuluJ/
lP9GeF0091O5N72BItWt/K5EWrmysSN/EkndhMFibPDqLJRvUqEQQZzPUo3Y67wR
oUSHRCZvsihkSCmN10/Aqm2w/bGRrGQzK6+JJLXSTcpVeMzmAiRDsIWXI9ZM2gCM
diPSfZlZYn2RYLxQ5E/864ACpSu29I8WWT6pQV7hV2s+sYxB+xyxozCTY6JSt+P8
X5y9JckUeTakF5O75C4O30x7Y23HTLGA/CM7Og9QQnpMa5d0v92X/60SxzrwafTw
sHijQQIqe/zTZhcplSlHnoTEq82QrxIDvfHr+pPjv9lCFI2SbhEqe8J/uyMRWpXf
ZYZ22oSYedpX50dTJ5cbDidfPZuD4ToyY8YmGUUBx4m2SbJcH2dvdjqu5SkXR3yw
GqmJVHKJHV8pL7aT0YCcOQwUnxjw0elldCWaJnEshQ7spXcHyCrR52WWItNAVxNa
NAFY8MITzamVr6IPWzslbCve4tfKf09SB8uh5NqYAsAsxQPP7Npee+aDpWtkbosq
Buh05VlTiXpvqjn9QNSn4nYubJjofchdU+rlenru1kKx94Dv+/IoRkTXK8BOBQ5I
3CdM+VpiD8iEvemumZduSdBV0hxqgoACa4Kpzuis/loAMFALFWmBkr3CjmJj73qP
5HZK4nYxHep3q2BUT2LCFcyXcG/oWoIRJ4dwLh1vYzXquILhWabEnbPwV/h5EM7g
kG1ELnzVz8IdC5zts4WsGJ9y/iiR1oczTSKqL4ALRVcRaHHsRZIEdrOPCYFHS1ZX
W3OD6sinfnZbsQApIo6TrYBxUH1n2pdIXjpC+Pge90UsX4FJ1aP79RTD7amKL4Fb
vIgWs7CDSlz0k+50GxdzwcBw1i16kquOLAMT3gU5ptcrNJCjazH6na8Sex2kwGrf
d+Tv2IWaDujxSAnV6I0wjroTRhEKR+wIkdiSaqmPiRY/Pv1vuPXLCv2fdEEVR21i
NFuBHHTZCmn81qanOO0C/JDesjhhnizqAJayTwcLusbewLNwr5eyegqvA9ulli0N
T/+UZEAT6U6d7UNC0D+SA/hNIZ6t5X0TwLAin3rlo61XjvvPmyPv/W0zkaIheE6e
d+kHk+64As2K8z7YUA0mCMNBisOfdS/De+6vLPFVH+tEHTgKoMwPaeahQd7T2kvU
qpliufvKtOhpIcdMj4vw8ZtNiYtY8jWpiTcWZkeOr2WB7JCerPew2rONvOKOcThm
EycBT71w4NsgVmala6CtErecL1aoAstnI5zmSjlPqBn35AKjZJzRQaMyyz/ynQoU
AKfTpKKfyRqpyPxWHCATTo+hGY7pPZ9uwhIhDSm1aPFEqrNkKmichaTpJdx1ORtd
wkzynC58BzvJbcSnI3wqZGI1csTAbFFD0I1+wXSNNRKxP7VU98rQ8Zet2g5i34zr
uLlqzzjD/U3wK2JF6vGbOY/qlA+6snHBMasA3fyqbE7fa606zYIRCv9PL1MDm1q8
zb3qjbP/ASn45u0pG+GjHSieujTUD9M7bN0o0r3D9GlYqNZjGKRGgOHGbw8dOqin
r2zzB5dzxStBEAXoqgvDos8KLvL/ZKpTR4tw8w05EBVSgR72CJkz8nTW5kbgs1T2
TsGLS8IH3/r9M1yLevQPqF4qNVmchyR0SH6U76TFxt6TIQtZwqt2uZN6LfDvFv5/
SF61dxj2NAyd5NMpYxc6ZFshPtRdAqC1vOIvfMUvXCgFfVahoyJ+3fj/7BEg7jSa
/yjdk0hBGcQyI2Al6z64bRwu7FAVqEZtkVx1HxvAIeyCVD2OJeawRgU01CjMQlxR
cBXbIIM3YaTdcljKjrFc3SIfcohjMZVrOSsupLseKDSDLrWuzdM0f16/lw/YIAdo
7rFOewjCTe5mvxHHdO3VaV434FCn2KH9VGf/m4MS/yx1c/RX7Nex/9TahyJMAH32
n8rBIvMqasxmFPLrgKEwq44/lhCzp1q4c+nyMjtgYgA/vOe3TkU9Dtt/jfbWiWL5
P+LrkanEf2V8BPhRwBdMadK5S3I2aY/l2k4I4TzhygcC/fBH+E06dd/RH9cRY9NG
dbKBz4DyOchaWoYmP+y+Tb11AQ34Aw6KhrtGqcGSbsVJLgsMMU2pyy5VneWG8s0R
ym9KcWC83v6NwxeKHCM3eJjAofIdUezLhWGvEVEq6vXiloUHtDbs33qz7wtC2m6e
Vv0ZkoD8yxousbWSYlK7oEcoSOW/BcRo5zKTCowU+2Jj7nfaklh/EAj+7iGYwIXS
SicfHm7WiILAxNZ8jwBqtIdcsGaxdOGtY/lpviX+QurK2q/8D5FifTIxFdzX6PBj
IVKSF8swH24MyuGrjiOHI1sTijLci/4NiwwYcOQwGMlrNQ6YX12udZ/ty5tUsnF5
kJ6KDEOBjOVbwIsXRDM1aOeL40EGl8mvHafxp3+NGg5DT+toRd3I42uqOlucR1Em
icH9mg3RGhTd5p+dVjRDQryV5ciCdcqYt0M7+XvclhMrG9J8go9RNItl+AOsk4cQ
HIzoCV4rOlqcmInMyvbF5WItXl/cZ/d3fTytTB5H3g7m0lo5eKDysmWsCXjsRrdv
dxktXs9q5/miz71BDO3tDLqmoI5EosnoM02v/0Kl3taH16cDhWgULkK1uNfAB1Bo
3Qin5VBYzqLFD9PUhZh9MMoNO3Z5fKQZNIoLAjK6msVsbJKqhkp0npKiGP+8N2ie
GthSdDDxQTXRrGIqTFzNIHbs8u6cMooxM+tWs0eIydkcM5zHe0T/uf8oncdwtoUH
FsbT603iorryZT1+PNT0zYk2u1H3flCPT9cuqwnhh1yVCHkNpC7bkiA0mOwIpMa3
OfOnEKiiS9Bj3rBRvXNeSwhZ1EhwlyixSiaEtwxRNvcUf2Co+j7mtPDLZLbO3CQZ
xynV+w91eKMW6Adummph4v2MmPN1JKriwMp3cNw8glNJZVsUeVs/wQ5jmVbQsAYN
+2H/0mYuM6U7picb95kUu+KsJJCKGKA3mAJqDHTTtie228Z1P0NCAqC2Pnk2Fj9s
07dLLIm+GoBjjirjWhN+Ss0Ig4CNQby2Bb6hUqohTAMt6HZyDGVdMLpSkhd/ykkK
q4y9Urd/6i/fi3BLNDBGq8Ci8e2qz3kEz0YDiBQE600glVWrH+ZmgupEJrE4HTJr
/vwD0pHL2B6O0c9Qju349CnR8ak9QOi5rq5sxKxdoSrxAG/Xmw11OEAUQLydP9V+
EEA/eiRjX1gnBAfoJAFKD3oQKh/eMq7p6INRCTFr1Z6esZ9XUXHiEwLq8z2+uSgS
M2IvvKNUxSqGj7v976kn+bkXKSGZm2H56j6/seekCMsvF8WoGjFUUkMgfBnNy5td
tZy0qP9QoWjc7SDKFSivzX4j0zPNPb7GOeFeJEgSwIrPJxKUokaQKUOk1f2p1siC
St8eDGrS+EBCtpB3diLuotQTlPqE2PuM1Q/hjmgFEWzOVWmfKyDKlvLkGaQ/3bkz
4EN5PQPd/ST5tSSTrs6/Yxpzx/1dA964Rc6Cn54rH8wVkZVp71R2BVkJJQl61Uoi
K5eVPj5o35ShRzn5q762rs8ji3P6FcQZidtaYmcLP4xIMuj/EckJqkvQKBZQcu00
nSUQbsjngqDQStd+WWG2sZY25+zHl5XtXQeGsKmp7j2P9xFz6//8rDE2Tkx+m/Ek
iHwrD0XE/m8PvdgKuvMOFEguEoojwOx9oQp/UyF1igUmqFfLNNmKNm+ieUswWb5B
UuD+06hDDn5lhpwGpcedQU2DwOvUga1QWpxcrP+wOssK2dFxCQd1BPODVp5lVGpX
dPgM0PrRvBkchPPjDcmpzbd0EB6UfPM80IfTxykCzxi35g1hZnrv8m/li7O7KFdc
pLSOckNpI0uU1ASEDRS6LxkGlCrZ4HNloMSoHvzqYEq0HHkS/g/1K7CvKiqlY3kG
KWNuuo9OVJ2J3gQDJkHevMqjCIy5KHJ9WnM4l9feQsFfqnCCK83ZiteoxeZY1gmY
L2GnjGqVjkF04a8peB540ox0wYgvU6JX9Wl2oxnuo3ll1/Y6DBRY2LxpggV+4758
ZeiIHdsF8MsdKnE+gqB3CAEYYtmqcbqS/yGaTtaWNV2cI+yUQ/k5OwSdlRvZRNli
U+mbcLQBW0QsnydixDSeYgGuFxrma+U1PyI8BLuMHZE+MF3qOPOwqupSlACPaFCF
wJdSIrajRIRChYL3TLct3nhGjzcsPA0ipeEVeUf1WJX8FjaInlWEcrLYLb8WJjO+
SKN40HEe0wn+MvJvrl24ETWmSNKM5UxyHFUqM2XDlOKmGXYiklzaWdBOUNMH7xyh
1eXec6EODm7AAUhrhNIFc/864Sh8IhWkBeFWo6/BnSAvH+txy6BDpnlO+oDqh1yT
0NzAVceI9GCbzO0E7OQMxgTFnYBtP2D+5mNOmn4+ce17ZNVZhRK8lDyxmS3+VnAH
HTRFDf1iCkYN19dCEepeMwEvbBSaDf4ryBvIuZp5x93rHA+DEvKg1DDWDlAh2xBW
XNyRksShWBM3E4bEdxQcSaiisdtl/X7T5DBjmzKcuP7I7l5sOOuqdwAoUjDI9RVX
zYDEolbVq9f9TvqJaycsAnVo19SxE1Gu7oiUQem+fhZ8V5fg2p2XcctJIv6Ui/Ud
Nj1DeFf84cRFTi8ycSDqhxsARDKgQ/rVR1nM+xMOXpk886sykKaWNQQmipM1ABqn
6aXWjMCGz/dgTj+sMc2rpRKYoS1ZFnf3SVvAFifY9VhKwSU8X3zJMSVjaii7kSf7
g3/kTdqIr6evSj96r3cLWsE+knh82jar5lOPbQyZNiUhjUJQ6pkxuizJuTgkcLXV
jtSr0tYByJUo0odw3Kqw4bfTBmtgkyY1EyHPyZD4NLe9JKR7R5pYv3LR4XGtjxQp
li0xhc2Yd3qzTTAYF956Xi7bSYHoNg4FMib7X673Q7It5K/W5ubZuzNZqTHe9cQ7
tdg+xYeBtuOmk9fW9OYiOZ5zDWdTK5TPcRaWKypR1n8kAqK91xu5LUy4Co+fT3vi
dwS4B+GLd8MR/48WYBb2QP/ErbhrSzi4aSUwzPOBzvRbsovtDl2im3xYoPTNcNVb
b8aGHy0AA4scRn/kpVGakwh695sq3Hc0rJca6FtXTt6P4lRXvWnvYVE9LHE6lOHX
0+azpxHpbCi4ocls/SayEzLXrG5d80Zw8EvNuWGYg7DqvOTvKkiswTNic+XiXkZR
ohbylPxGwo6EzB6KWW80w996ckzDhY+0KyCoTTnQs6ID1psxEhqYj+0dT1SmWMXR
73bGqZlaYIZE9C8sNYp4T7tIUNm7uuXzfQlTxd7t3+wnJN9zuEoJnxlDOoMHg6NH
/YB4Vl9uvtvEjcptKWc9a+A55rAQyKHol1Q+Uk1GpuW0LVrShFX63bYOKwiN7xQl
D1CQZgwhWbVjFmM4WOaCFDkfnruSP1iC61e8q/aySDh2FWztgxpZueL+OWaQuJtw
TmNqSXM4bahpfs0Cfr4RjSuIW3S3KZyzuPyOmXKqA7p8cPzGT4kqmY/tunHWIpjs
4XLO0TmkM/0nNTXBB+G4QKY2v3aQUHMo/1NljY0AJeu1kBngTx20beI2DiskUd5z
D2GwJUOiAB1SQcCyOa8TUWTFK0LRnLbzaZ6kAi2nHn5AGE95i3XwEyfGj7yT9ysv
XDJr/hdKzOwj/uDvKPJOO5pJ1nlO2fAiYbvStecAdVGfJDXj5TH0/m7C8jTpaClV
aiKZMgdyTz/wmrDtXwHAae3cu2s6lhpIFyiXV+7zE+5sO7uq+D70g07EwT11guAG
Um2fKWqI5rUyFAbb8hHjAPGPaLNAawL6HUywWIyc7paIbpmSpyMREB+KrFgRnkA7
YzdHfGjY78DfMS4WEdE+k/K+07vbCCBjbfdhBWX2KI/5QZq4uz6kFGfvDP+Yc7h+
sAsnBoXX/wlpmw7PO0IXs8esg7pvCTfkl7WlJJvUNrCYAO/siWf2CB2b+iANCmRh
Mg/q4MG9aVvTrS4NnqtMes67KVgCuWu1c8cdmBWHsP4DJPb2/Fs3x5sARaTaPsjG
z/h6xCuYGMB4dN1vfSsR/qpFgIvv8mPQT3L+4rr7cTbkp6jOi8L8husCbjIi08pw
6nc4mgsEDkIwTXVqEdXiK6DDd8ZItWmYxUXfpSafzRIRP2V0lPPSzUp1ImkQNNgT
wY2pwTfRlATLMJwElD/rxkJmKiWxy1Qf/SEpkfK0f9SybtXv5SPFAgtyg9aFfbSZ
j+2hRj+Y0UwHNhHcCUjhGhRYXzEF8ZN369piSqTnG30SWYUpcthIjC5JzqsQt6GE
WUk/6SdahZfjvAv7T14CNyHIDF9cF7tgu5hSBBRwv3TDySW18523a6ytxriQDvlh
OhzIm44qhpzFL7qcGR/KG2aUJo6SxrQAfpRlH7RwH2lw4F2hEKzQAl+6mXL2jKEX
IIMUoUOVsPkno1pFdvZRABq3BUCxsApogvgJP/bZMfpCpcbFe9z+pFz3L4eQWXR6
CcFk8OHf5XfFuJeaiJvEF/DR6+qWGIWn9oHEJP1Reapv39vKQkZUSlUpC6jGtnFx
zI022F0ZYL3EU0cHSZNBdXECUx18daVSsLSsnXyXeaFKQ3NmuVYzHBMoY5mXW2Dr
ShRu9+n4BjLTfwTU+mwhFgBQkOiiz3VROhVoH09bfXId2faCGffgvKfwNVfARsJw
FK7QtMUQpAb1RGEQN1/rvZd07r2OG6V0ZE/ExrOfwFNvdGzHUmT7UbbadeiksHHa
+RRGqyhIXoWeFuyHtVKvyZzriejTmYttlk0fRltop5GXpzUJLV3AChtyQKRL5c22
5IVk6cX35eGko6FplK1hdKyd9JF3Iv1zCHDQPGgj7Tl6GtDQfdLNy+Husz4dVMls
AssSZRxGl5pBMl+OCFXk0KYi9Ge86mROaU738ClroiEPR8RUysSz8y4L0iK/Pk3o
KmdD3sMN4ZTE3/5waf4BBRg8P1ZCNEnC+TCbYb9DVndEU7gLjOgajSxDOCmGordX
xr/o51qAJYOd8Q9v3YYPElXDiKU4qvGAyh1N9nLZcnbYVFpB3Yw868Q6IFFw/uOW
Uo96AIOJRuQXsY1KX461JsyuZRaSql8WMaEKr9UHsDSBk2ha4HhiP9i7UfYtyF3Y
5xiiig8VaP/WNb7e7WsiavFtPapjNkL1ikvj/9iAfgfHGKtkJaVRl/8QUaaMJTBs
X/Y9FNUgESaArgnHfWJZGC45P64jRUe5g5l5kCSO1B420UJn06ROspPXlBvK4C6z
ZQEzgD/eO1O4dFlY5plq4RBSC5mx61mJv1F/aVJkWyIE2EmwI3WT2/GyA4x4+Q41
pwka7ySphZljT1M1AXx7FAi2z+iGEB0Gw2yrMS7hlnCbS/o4kqmuapxQWX8I++Gx
UZx9zJb1kKHkvQPJ4tFHbwDF5ois8KQRLPnc9citdCm1dBI3/Ro14ETKd2Faqd7j
OgCehCQZNnYu7RONVSj0QsbT8DBJMWrdTkuoEcFloCFWrgHTSA69vr7F5NaIl4V7
cPHQpZmxsNjjuVhqEZEAxr3woiXdlP7Hr4Yh4fv/pO+mmUFdLP7MDl0fv4kafMyp
V1aVs9hOly6bxLb3tAI5Oja0MvrQCc5vt6/oYh/83AwjYLCwLMlp4RemWkEuOpcR
834V7y234dQNBy0AqwBBrdUDITEIrPNRFnRmkJ2PvDgG5d70FKjr7at30BM7gG9n
+s+tcW+XTDbgu2Eso564WeLupAyPEg+Z6YD2pQYW64zCNJFQA19xWa8OuDd2U3bB
DzP8pko9Z4Vu6WyXTb9HXkEuPoc96jV7NHNfeQdX8tmfpsFenGgEtazSTWEUEgXC
d01r1SD65RNmKHKOkimRy8VdXzTAri3wDrKmdnuH2qQToiLDHtEp0i4oqoSqlLmn
+MZMj5at0Tp4flOT9IFhviwYV0z324pJykNDIxRBO5c/VRXiBiEdGfuxcKLzr67z
YEFRAx4mfdLMxpcHDuDz85/yzCrsdi4x3b+7/XNl00OwBzZzq1ZYoLpIors+uTZb
rbwO1C9Sm+j2F9A4J8sAwVeILEbNeL1rXDrlMWGrjogJaNVncB33sord2zsmwhTW
pnum7k2S8KC+GndtD8kpWya1rmxrhWW5JzpW7pP4aSXaroPMk2rQpuCQdnozUyw3
B6D1uh9H0yCKoPhQ9NThtBnCJgzhMU4D3vIUCv6YqtnNqOED++zo4YQ47OpsYc61
FlEwlkR8bXwhd1wR0v3S5Si+jddACHjFbg+/Fes0dfvW/acQmuaZsfkxbOrgSmPs
dByMKHHU3/Jfdgahv4RHtLDPzLpfPbhUn2h9UheQRZyIwUoFUQkdWUltyBs9aXil
RxIy9menk5u9ICVmlCc49kAWl4qYlW+cPg2p6BOqAUo+isoTf6IXWFg2N+TJXk7/
2fAT8FFDKnZUcQZ0FnOXQ5fzFKGByzKaEZzkzBlKILzKFjXPi5NNH2YhacSNVGoM
aU1h7qB8ttZSYm/2TYCHWkVcYXfLtzZwIUXQmHRYw36GlJfmFjQ+L0JhA4BDvQhG
uU2B+xYTBVgBP0R6gdS28xWG0Nt1Odp92E7mZPNGXpTgaM7feu6JND8rtoIDj87j
ZypQPKgcbo9pQEUCDE1ZR4Al2lRTIjgDgbz65j5HYDZKzMlCFCk9ajdlatLSs3TQ
0h3xrSOkI4c8J1EWKi6nGuHUUtorZTLr7PaHmddP+07xVZxHC6a4CHwAVXADYQjE
hwOQ+fNzFJp3rLg6exMmXjA/pbh/tJo4u7BygApwSNy+k3KTAWDym6GHBqQVqXt9
93VLXbbgB1AeKXhXdVWg5tIJO0LR4eHN3H4DMDRne5zB3vlWX/7xr3sO3TW526J5
XLuUwjGICaOIRRC32J7AR17+IfHuVvxDWxrcC1IZN/tzsNcwSF909FIvIrphsN4y
WrU3n24mC75Vcd7hlHLQmMEcetseDFaTzKh7a3rDoVS+rMEKIBZZfzpAnvFjeGh3
jkJSlgfwHBaG4eEYMobmNehMNIStuxX6PDO+gHETtiGInH4tK+wE9dFDArFz88Y7
+5ixR3TKMqjRJoXCin+iYHYFHvHqN+vpm5SjKUWVEGdUTILN0JqqLKU0GzxfGQdq
fbl4z5dsipZ3X6TVvq0WTum9duY+SnOo8Lrutb5LcXVVoYxybKgy6BXc35rR09Ia
v3jebHUeSC+//yaRhW43O1l37ztFCIqR/MC2mTvYaouofnTnAJY5kQ0sk3l6h7OZ
m+jtGxYAPIPlpzDgUGcio2TDvZ9k1YzOwjT4piNNdem+ck8MOuIc2ppu9LndV8cx
4uu2R9Fo+YgzwoETcRR1AJg7PjyUMYSgr0ljqjP8xsPjbACDuFXpuu8EvspKtvBH
/9QderaanmXB5oWsCIg9bXWzz8dRESuP5g40PdOwwSDOBO6ofu5ThRQBLHOM38zk
G3TRPzBk29JnkA0jSXP3sYM0l0+eJMszGjtrsqMV+KQJOJGsTARGSzGnfj+oV6Et
I2QGcJTdal/JbJjEjGiQmVeZ6V9+v/s2lcR3+3KRvx7leYjLXUlE2JiLHlgb9c58
ezoiPHiKJJBfu6qtX/tdOcEPiGp4k4gBEq1dH/jLvb492+uF0R1AlxL42JESt39c
U5Ay+rFsxQIS7y6FPJoxWLX3BwDZ4riG7NYDH5RWwcaN7PskgYexSOnPZyln920b
uPeRtYPAmZW/6GLYKJig7mIg6/07k51PWEP8X31/pluNa4HYMXEeabyYvI6Y/mWW
AhO8UUD43riwZYlBh9pmTRO8eXa8L0/1kvfPvrmst/t0GlsbggWuYaUYI/ytFie4
IVCpwCJP6/xoszsqNcXedGA/h3IEMwexRiXNbGeSGbTAMi74X9Z+XVbK4T6Veb+0
FO9y1hQDqrAeBjeOGkAu32MrSg7jQu0X3vXmc4Z90k27IavQKkrUU04PQgNBR4Nh
OLVk8VofBz/8TSOI5hHJk979cy/CVwd1GrDUE6O2ozTkhE5EQyhhDm8IIxBla1Nd
k410c07G+IGQyOuguIgbDLTUGrJ4twwim6MxigkpfoMTELmKmURoe6bFS+TxddpO
kdo8YJwWSIC/DD2jaSqA6Dwox7Pxlh2c+0xwCFNCdu4CI8LkzNSzqofXxiSqDW7b
eNV+6ep1gVKhSI7W3MSEGfZmRZNfadtRkQU2o3IWktCVPXEtPVa14H/UvWOqgrUq
hFnyBmVr0NM77xsfVU0G4n26i1doRDRYtLbLHDeuWGFXcdi840rjlW9JNnJLuSHj
Wfn4lq2/PgZZ4sPj9CkUwJq8PURfZAkwxPW2SWkGEfYN/eeO7soSBeWTuktt9JZ2
91V7sP/cwkqVBcUfJV5S7hVZnW2IKRDLSSGcdR9OkH5I3+NtxJHEeIXA/atFNpIi
xqbbIFTZU2Lo0uLi9DvaONAG/gsRVotB/DyUWnY441q+2fTX+RayzrbsYUgcJdji
RrYCcWidkB6JVHUtMA1vh9ixz1pE0rW2nHmj9hRAq1o8xbHDNT+0lGqWJpLUpvGp
wlGFTx4Ld7+mAsKXEzLFGpLak52RqYE0Ul/2WUO0KM4oVu/5ijVSUWufwLhkL7II
SZJe1wOrh7BiTW45i87qrIsfxK+0DCyL76akYCZAbJoXQ6TasktHu0tgJSg/14na
nkpLkNT62mf/EJTYV1+Y742jYycgP47NK2Njaoq6SAZOeB1IfS33EXOW8pvSl6Am
Zm7HPofbO8Mh7uXVSHKx7hQwehUrA9hxW/9pyfZD6wMV6S5GnIG5oBPEJ8LADi+k
koOrKQLz5uLW55pepO4vppKgqCCT7lqD2JLIwuuTqZ4HqMXASp7w7bnR229CB16M
6BJkgtsJYK3xjohSRL/Axs9oQXZDBuQnVXqZW3OaKDYIzHncgVE2szy7FOWGeKVM
ao/UY8mC9W7wFLFH1wyhnvQD/iRTWoSH7nWw1bjpL6YTuvEoRxcS+vqgNRHxltHQ
rBWeuF4eYt3GUHdiQK8+BLWvHjvvLgr5xh8Wp1GtF8gFkz2dAIf7oHLYsgsT/ZHs
c03o1qm+eO4KkMMdkGML8nDw7fB+a5wByQ9EnHClLiBpx/lkSvYYQCcq9usNpDi4
EdNJQrzddfLKmjJu7b26Ah3n7uiD3oamdPc3g0jLC1D4TrPFXgLwwYY5VR7wa8ot
bkAmdpqZpL6D9E1GlVxxX4UBgWk2zZ3HC4gXKOlsL4yUYeUxcezPOoXBO7eNaJil
OXDa+9otGygejIXJEXPz2SH5nvGlRgfHPoqicUrVcMipadEweoo/RzTfDrBQWVMd
Nqq8M1/tiFK6gHN5cUvv/gNSsU97C/21jZKP52XFbSzkuYc4XdGA+T5QUbDIja/2
O4kitx23mc8ub6JJHp0QmmVh6VEUybkv2A5Rd5nkOPI3idwdONQ5c+X0Bd7wbd/J
9CES8fSZSqlqbfuIPiFZD+TmGDByivDZXBofcv/6BK7w2UNYqJ2zOcN5x7DwCG8D
OoNc03UVjTYf4OGbF5NuLsXtoDEugyvv6KkOeI3foFE/SDa5Wj07Ii9fQv3naxDf
UDhwcXL12fXCK17gwjhC2pyemBUQEtKPVOzAtBFVXXSakTU3XmPK+XNxeQqYEUs8
L7ICyqxxH48wWnwjj8R+gqjopi0feyMohHU2RPAbrTBUKmdKuDKIwBJoGV8SVct8
LH0uHmnmJ3b57yPH8FVVXS9Rbx3/0BIS45NIKYSJGoBC1lRw2m8x7XtE2xD8QMZd
/8mNUYrYa9yNun11Y2U5GG4cw2dVsdnSqjdFCKMCrf8pSVjqJ7lLMHN+VWHQb13p
WTIv0ucwJ0yb05n1YpwC4vHxp4dk4NYrZdZQ/XQ4XA98NAXWtOQvroOLnnoJHwhB
t8ciw0aY7FvWzUcZr+LbUxyAa41+VKP96YGGvpzCDBF79eh/1wQh33igYajCvjv1
NmueAAt5bX2k7zs7axvquXdOwHw1VMwlxR9jx+cKKfaCttUDGD6CK7bpSJQQUBQ6
W7v6fCvRMdcJMhudngXkZcY+7//MQncIn3x3NqQ6mSv4vIuehzdXBbK9Uad/kxLq
Z08Q9RvSAN3BpW8Kr8lE20G8nSc8XEoru1BLsoks8RthaOmuIZBHTuRAkiuRSwrA
6523dT/Axwlyd/HADqcwC2qblxlZDbWmVqcb42JWbRqi/OWF3yz8y4Fc2mPbyDCY
oizr1GpXauppv71SSGdwJpWsCrt48hyxXre0hJ25pDnH/wF4IX/6XuoIcjc30JVg
kqWQv09RpWbL5hUDMUesJxV5w8WkvDaBis+0wrsWNBcDbxVDAzRB6ZLafjE9sUQJ
prXwCA4c5a+A+D2EJy8qHlV3/FPvnIgEhIY7R54vnm/qNLH21Veg152Ggmz28oOn
V6AEdqSLYfpe3IScxOd1XOlkXJ0EgHZDk9ZSBWoVKS45zPgQ5q4usiRXUiO4pKLs
GTxfGuErJcsu7GFt96v6w1GQ+mx4/MAhaQdcyUoMf2KlCZ12r6iYa98Feh2s4Sr0
ww5PF7iWYUOKaWg0BYv1M5o6dP11HtSQa5ntPnjO1VRxvgmP/pzJPtZlKMIGWnxw
hGULqbGvavrmcc8QLzFIhiHzrF5Gniq1SLvL+Eenf2mJQrOU16+Ylv0ksoI9EQE+
6qe4XRVZHXFJuHBhPf+2t4mJZPLD3corMaLInzrYVa0lhKqtrSudqEnGUA4sliDg
1yVTndZK5YKPDUuu0ANluJ6szEJ/PvnfJEvBztZXx9fT2U2fi8kRHle8XDxKuDT0
8px1bQNhUD9292OVONjp27ZqUZubS33v91Ow1/YL0ZZqAzl534Oxh24cTAJetz8u
AdNGoEij7Hltts2Q066WZj/b/eAPzwY+1cIfrzvRHCRPbaKNG2mH03ccYivFDzsg
Wjz3Vk1DI1yegs0vA+ckQF2MLiZ3Fi6VrvBO5oFzCOBIokTgZwsJqINyO6mUvbK0
JkVv5bn9XqwbDexuAOWU6FqXyL0XTspJMlh/iDoiArgbhXEM6WOt/oMOkMirfMpm
V33wUKAlk5o+BZ5Khc0OqjaYjCPgtgIn14KUuvCq0PZ9TMKBodNpY9pkjef5q5rR
c/ct9SlK6n3in7tGt4lxxS7bhgopNr9stQiSttyQydOEth/6THEPvM7I92S9QusI
vI++3s/kLqshqvHdt0lwcnFG0sme0HqMrSK2yzzRPJFkYjtoaMx8Dis6caKor+5W
Y+RyfCUp0dvywh9ttC7ariuZe9yDsG4/4NO8A3zM/IAB/v55lfgLuCA9KNc1iIpx
4/+PC3X3P2X8mpDH1h1sGPD01hcuL0+Rt+dOAVf6cv71mUjrPro3WRzYf16F4GPb
oiFGu7o0QM9/fCjLcnFAGk2UKeT9oPF1fLMe5puK+9Rmcbwt2ri9HTSTlO4u+9Ni
H9+dQBevE9os1ndO4HTVc3elnYTWb6Exqa84DatSlmG84RdCSQHBJqMZ6JFfXe3e
7l/k1kp90jMKXB0mmXEbkPSqKFS1UG5oLTXGdcyLf1aOkTcnERjrj4GnPuF0ICKF
ky1IIElmLAelt2GF2m/rJYkuPfnpdWCceonU4FvvuK/nIIGZNJghWYbBWxSoMxZg
LpNQ0LMHTT82TMDfsDYj1fMoMFr01vMGCRgS9AIcG8lAKs1i+wQYkyW5K2D+tSF7
GhK9cjxzXPtb4rxfoHmpuHF13c5KLBn2L2L3B/rFjoNuAfPrTMROY8qNf8WXkzZu
3TEDs2sx4ZXldLkp2JUucP33k9678TdKkpfzN7M29SEF0djN8ttj467fc+GI9grP
ZmfC+rUK1eNAGvU4lkw56AHZGbg1mV+GTA6rMFu0TiS+8ALa8qJ+uI16SP76PHbz
ImRhxi2LDG04Cwgc423xsG95HdCtr2edbkdKbKuas8FPr+O+GfYn7nzkWTU1LJuA
312XcL8IZKItG2D67HMoBF3oYOzG2cqiPTuH1sQzHlbanm79Iy8LBysX+D4Imw3x
E7kulv4AtrGA0ko4WOaogxuYjecRheJZjfnevLY6mUORLLP4Eoj3kkJphiGBkGyg
z9A1kjneWLZEhqXfu3SmCu2pt2PO/j9XoYUS2CdS/zTTvcX2OjVAmOZf/lvwcTOb
vZnbADyRds99fF2MOwTW3h1jbBK6EoffiCZqK0HP3qTIWQQxdVFYEyH4DhRpX0yJ
pfPrhzD+0jt83nLyxMfh05ZuZB6suYOBfVgspXyDfn0VhTnT6NlRNbvFHWS7TmuL
PYGf60/mWqBOrfozK6wxoiC8PElqpppvDnYsvlrEkRKJJckYBZRskmyNvfmyXu2L
lje+OKyE9UBwcbtHtCAgjk03stjNZdhfWNwfbXZRpl4Xw69cS7n2XbFNGA/xDDYS
lbi+5QdTfGbjphlhPE2KOv9rd9PO1tZs+ePN8KRe/cpgD0RFs2Udx4u1quoKrTnl
DUUvMqGtSsOU7K6zL81uBjappFLxLT8DxX7KUeQOCHfL6uTuezem+gDbgMxuim5P
JJ0JTlNkDv97R3jiUbrvhxiCFY2Sb5S6xWNmALwnJjyaBmQbboWaZmO/Mqk+zZr0
fuCyMNPXGLtPPANeU9xJ7Z7vfE+QYaWJdKdka4EGPpuZoKfww7WdeWFsBiwIFeIb
2dLSgrKqdzhlrqLhEy8lEL4dAO6d+5p669Lgf4vo78JRImt/Kglo90utz4bbSgpU
nWcY3MRUHYW+W1Hhk/+VD/fX396Hfs1wFsbI8vQZyQHls6/MwjrDeWs9mrA2sFSn
3IRG/ed+YHTU+CZgEs3zeDrh0d6Ubb1wZeT/Hqowcg+nrbDarvzgyfD6Vnixd37F
StXEOYkLJvjYvKX55GfmxmxtkuaCVSiZKiTju1rjQlBsIqd4l+DV9BI7fyHBAHQB
tymT8vMDtMmLsmlyrueonUDgWdyQ4yJEX+ogEyqHqqcJR1MivxQlYdmoRyG09qA5
hQVAT19i93nPqFskdVv2x67YlXQKRK537oJjQ6928ExbSfKmXuqdwaalc8PLEMQU
XsoHNF1A3Ui/epCcu2lrupetX0b+FySH56R51IN1UFUjDMCx4rnvMiaGJ242f48W
Jtf6ZAFvp8AvGmA4/T/YUMir6nEbNLolwMlGQdkyTurYGhrocpummORu/QDyB59W
yUDDDBc/1ROFm4/UkcNc7p/sX1p/n5XtAj7/e2QGCbc/TvFDE5xwf3USKOkyZRrn
Zysz/YO1vFQI6jvyORw7KvD4O9n4ltUg6bxK19Asa1q+dr5IdNUUL2vFDjhetOkx
fqWshwqX2SWs6qTz8rYug1Qm34Qyp4iI939GDKcTj0+NEU5o3Wx9cfGXWjG9k/Pe
WHAYJwileA84oO0fF5IOMrlCppRnzE98zcRpJhn2YDSAorBpPpmfNQCO/wwBf7s8
4xiVvxF0I6fPLZTGsJb+sCgdRQjZi0YsGQxXh+aorKxESAI+w8P3MBHSE+x7heGh
ObhksqNbf6FSnPE4SKEUiY5ekwcW2raJbtvPpdy8FvdqF/EQAA8b6hy+ccHagOEG
ffnDNunO2YE3cjbYFR98JsSwuccjBMGSXgph1+xoa0DTMSJIt15IBJfu0rOjoYuE
Jm5nMT5iu4dqi1JdgYjsrRHo5J8UPsSzGqf1imxwYrK1i1fK1WgMt8dVZGAVvdUd
dGePzQ1v2Q8bTuaSedSJjnngYahg6Z5lzzq5AynY9yY7A/6MQfoTYVQzFROrbToS
cBiJPXbW10Vg4LcEZ33oXXbDTXWuYHVzdSmTNfxjOkAvcopme94ph9tlnN8ehxYi
jAfwDifUZCAPjUA+3Opx9y3raA/OiKrqdtjXFVwTHZzDzT1PbyzMPnW0JrW2Fktl
CkMmxQhQDvB/EalKVmzgMK9eAhrc+sVWMSnxndfmk3LEcxGAesnk/VpTGHs3mAmI
z5rNBFzGZPQL3UdRtFDcYD8osS6tlPgFB/pqVUC/DURJl7MwJIva6NYU/YrBKln7
NTCW0J/jNuWDSKwPgXNbAosGAd2gXrH8PjXKuNImoiFgJWkPQeV/6kKbSwmZ8a65
QvaIAEvarsb2hjhaRmTxeDOeQRVAmiH7xyfgekucYVdVbmdp9SqN+lnfOWF8GqMr
uLq7lzAc/JrpRzbvfCL0zLPVfllXGlKBsPCsQ2slrsbInALBb92PDSaSZvq0CuLU
TRJWnB1336LcwXs1Ndf/hltLVIuP8Kh78uRkvJyeCu6lpvorpL1wlCkV1D8WSwC3
TY9VhmRNH4Ga0xHB/7okklG3W40JKBw33VDNdQBWasGTh4j8534Ae1ylyzxEJzHC
+XSk4BI8vFGJ70uOCl51/MScMFt/K5pOrqWzvLIclBcpwcUVx9QWQviV4Q/2kRf8
s8l0LvjuhNYd0sBhsncCDEOlJTBYECO2os51+MDf71N0L9b+sLG9xSzLThUTMLW7
CV41EpHMnDIEDvwIKcn6rSmHeWiIBBspQIWhzvZ/KdktE7L4rhzXe84hftTQ7OC1
m2iUPCMjEjMq1tS3cmHkKbAVuNUviqzDAFnS9lum+boILP8GAOeDM3hUPQ07ZzVH
VUpURxupZk4LhGGFHtor64UTk57QczaFVPAY9s/djzbislpZrX/oC6DHedpTCzAJ
I5zvHlSJ3Q/UJBp773u1LTcv0YaBAl4NpbwOQXRxm80HrMzUHe7XCp8lidQr9wbP
fsDcLXz/wXTLd6XDN+9dAu4pYgTRgtRjVWQkjHlinkVPffambOIaea79xV0q/+pv
u6+EqC+FxWjndgOggmNokLy0NZHrNqrCCrOVBLsWu+o+K7jZyinq3hVgtmQTMnHr
OEI5nvp7VF1yqnOo1aKxrgta5wehiuspj4Fap8LWNP/N20OPeAyFzCbrNXEUZt+x
tl+YeCWLkMupgYgmOCBCQa1Df/XMoG/mC9vuRBBlpqm297psm83qpWxfmkgSuv9C
4k0NLQK5Wki2sgZg71bmy/UDHjOPv/1FEIqm8rIoVDt7Bil0lap0o95htKyEQGOo
ywXHfjJF41m3xOKgnS5O78cptYAb8T5dk2ZATlycU/uRSPruxuwtTKhJhwVChwuK
Gg5/9M3enQ/s6v/l0ttkwZWU8PUe4NRrEMlrAjlRBSsOps9GYhT9xJm7d/vHhSTC
PDAFmEr6wNknrr/jkaXK1BzaX759FaZqpJEZ5f926ylhoQ4BD9O0glr93d/Mznek
moWvVbcoPnCtqs19qjWaa98Wvtw6P2vuVjmQyo1oZ73H0HawOxNrEZJk+xRp+Hsf
3DfNNTkmJ4S400ABATkHNLlsaJMa1O3oXiYX5reLU6g+BrvLxm4LVttDh6CfHl8h
Ex7j5pzWLGhS9hHVo61yP8+ifCQNBUVGvTtEDDhfloM1Z4zvJVCaXjlbV0+LeGAJ
tjXN3hF6GY+aT+C5B7BPWyFd5WiSdenHxWNHeYgpafylRPKf6x3MyHQ9dtsTRzN+
t8Ufo8fY3HKq21cSYnNMlBy5IQn6QghCfGAPfq39W4cypN36a7kVS+AwjCoLpAVs
cVPfqsSncMYCAkroSO9IewTfMaKHPkJFj7WMvx/C2g3sRczbJWkyDbnA4QJRth8u
XKzC4LGYboUPypzjuWP/oy5W6YVRvLMoTk3/I3HCJsOnUaBy+QtTZtPJeARsoKIU
Y6WT8Z3mzaC95e0NxtfQz8qT2LSBdg1YXJiA8QGWB+2udZfIISqnWFWfkajOME45
N7YPM8H6TY+ocuakwIWkYqOV8rm9WZeWx+U0GsZ+fQbwZq1OfXQ6K/RJZ651OWGa
VURdcVnOjqqSWEv6w2cP4/5Ehe7sYI7C2JjYZEgu3AvfueOZCn7DWXA+WEBk+coD
yMEmb/883Q7PjeiRmCLLimC56rcN1S8Uch65Bf1uqvV7tkfkPENLNIYS2ipD2sjL
a1YDOfYgZQde/JLItfEe4GX7BfHVKxEeYzt5d+bOBZLgCmyum3pEjKLAZ48j5C9O
Uo3UJDsNDS5bPxXLhqUyhJcwXTHGg0Jm08RDLyOUWREtuos39U6Fuzg9ykmzRKC3
7feiFR0rAhIiphjRV/595ZNIeYp2NXyywbXrw87o8kXbLCHnYGJnbOYG+ZgYswMP
HDtLtffzGNCBupuSkARaU7l9FPscXjsEiOUGE1CLnIRhVYam7VRoO/XLzaj2h0pd
f7SGEWe2cwrZEkJTQdmNAPjlE6OFWC8zabV2GsCmKADlFSnXKd2ecxGNoJAEK8zW
UUKrHwF7PgGd505mcwc0T8NCzW9aGd8RDE5/DOaByGIXxFX647ej8Y1baO4d8OD4
E0SaWohZAze+zK2i5N/LkHTyC7/6cgW3RTqH43mDsy9b9mwG6HdxibMxBU1cLJ4o
IWx9TAgo6Lt2bjkPKEeuCxlF0R78KNVxkNQFuqkdxHP99o8dLj3ju5LiRFL80FhN
4l7TZwU6KrNOYVARk0QnqFEwl/cHzP+fJ6k081b50FlL2P0F8ck6Jy1wEdB5Ody4
Yzt0inqhbvsG/ajd/LUdMYJxnWFZjYif4mfXWq9gfIefimtk7nLYlAR22lJH9aHp
WZycubeLvNcd8bUgC0hW4JZ6JtXEY8EXFO+pB+5BM3nF25bRN2cNfDCP6Wn/Z8xX
uj6ScJRfNX6qAet18kgT811Lrn5eClidmhrQODUs23EQTcSHY2rYVjuOzkN2ry0J
IuKf1aa3tn8gQAamVgscB7AjfrasmVh89nChuknkynIpxT+xemDNQENPCyAUsRye
SRH1vitvnfVr60Zpy6uzC/08E8qESYABvf7bTKKv8Qlje79L8rQu8vKGl/HPGeYC
ik9v0BrUTePZ5GIH752lVrvP9ggreGu50F+JiLNdWLB4P/y94U/NJg52Yc8C7k5w
Mn+bRtzU7j4lDQ1ccKwDvxAB+EjOIwaYLMCkeSjYooDQtYGNKU6Q4GtCs9AFBFq/
hifhCVb6LttBeQV5GZWpLpiFj6eMf68VvguOzMok/aRXINR33RtLmEweeaFmqA3F
kiUXtrj+8heb/VjxTMLtE1vb4K9sHaJ0TJLRkGRy0MthT1qPZFSN2KfqBGVPAoLd
31Yy9IPuqh+1npV4muT745sAPi97fkQzU9pxRumk108O1bnBHlwdcetIB0uq0QYd
hsIBdTZTu2oArj6nr2APAL+4yQUvprZuXWmqVsvVJIRID1dEZIELv5o6q/3NcVHP
R7M4PtEN8MsuDOwdI2GDD3v1Of6gPU7TwrpraD/EtAb3O/0Hr5INzcYMufWT9tBC
2vfH2RZbi+7Ylfx/SKtCbDc5LLkrAm1cy083RcwboHlgLK27EexPfipYtL28I22v
RXp86gyaxDIM+XcIB0aiHfiulc2s1Rs2o5O+GBSleM1n7Wru63Dc4mfFuJdODiX+
XkIs0ktR+KJwzi+HXX5+mpJaFMc/oiIOOlIyURKjlk/qEQA1cGTNjWNJG8S8lWxJ
g40tloGxqzobc+wwgdcueItoCBH71gJCgYU0ROdn++IIjtQxbDSDnUzlSlH5Ib+4
9aIWSgpkIPbd1KbZsWZOuWcW56dxD9vUypd3vCrH+7e+miXhHxD+BbQkYgbyH6HY
0Y/d1o5m/pdQEkmmLZ9ks/OOOrT5UHXI463GDK5Zso5lDbKFce9eIQFPuYiITrHa
3UB1tX/ZX/jesTi7jJE7H2E9+E9q7JsODMaxQgxN+ZPAnmuRkGW3bHFTrSrKuaCK
l0Rsqx5hqUj2YDnQpi6QeO06y3p+fsWX8YQBS/QQrW4NC1PuMR8th/VtZSJZz7cT
nAvGIHAM/rJDxuCNl8VWi6su/wZfmBhbpnnCIiQqQqknJhgnNWmbKoNgzJd9amHk
w7Hs0xAsnHLOU4k38A349xuKdI3wXO2EIu3SmprB12s3UiwJZzM79l40R0Na6eQP
xE8eyPFtie3y6LbrEavFdiQKdcK357f4uz8VMKO0A0SsXcB8Ma8CIHdQPYpE5gst
lBtQswKjzg0+HIee+ZHhIw7qGbo0Hgb2njqDEacAeUBvslikoWZT88HPbBVI6Mpy
nTyCCE5zsDSxC3JkU4ZNGwPJi5W5AHVnIfB//u7q8H6bdLOQkEQsNNHk6IIw9VxO
+hifRsog6QjDRDxkLhRY0NpB6E1It3608ecTdae3IlLeoKwGBJ3Codf0YgDhWYqy
jQEasCxf0xFxIypjpHaWIOQsjYp+eeaTmWUnj4amoVJtt0gX0cHVNgcTItcV3wPW
EL0HSfJTVuGE71WtKMflMap3mc5piW0XVPIsRqBgN/ktaYjpNtC9qKjuR0UxER58
tgp2IntPilO6zmTygJB3sGbHtWBSzMV8CNeJRJPA6BKOtbtBuiHP2wegWKKQZojd
H3TpKqvYY6f/64t1IbNAmNo0lkikseeblUPq9WbiLTpJC7sdhWWGZSHx2Vih+V7d
C29oHd4m2BLpr2p3julRYm88mcOWxCYGiVVGIO1+ge0nO4UcXf0BPPeM+YpO46ZL
m8ht43uDRm2Z0UViHDTOQKF2WdCeYxKox39I6rcZbboxf1Lt6Y23ZhaM89AOt3qx
Tpz8f12/QbncPw9lFHQogrWdB+rc27DbKCf0v43NyndjhDEtkEbVlQ1IgGcI1L/d
w+sWy7+XBGEkAEb4+BQwfQmLwDPv1KqkLXYgJjo3QfMTdYpNeeV0OrSSvUEaGF1M
sNQZ1606kozbb0eDco8DLmOUrBCnBSR2iWEKqkDIjk8O5eBzsHvcknLdHnJX3+/X
2oO/jHn8o96lQVRbNI652hQQYnHxs8z4uciE77jt/hFpC6iYz8TCCGogf8wLnD9E
//Y6B4RCj7qCgpsFhtYNSvVIVHRmzZ0eURBM4SULfkk9fkY4r8KyQT+6ojJ0AYXD
wHGX5tljMbY6psBGbE+bStISWbRDpYdUSGtob+mDTyfdUq3inA9xeWQ/mQmb4N1b
01OD2b9A2iLkuL9aGcn/wT9UtcxFLeuBYNU7cQSE4RUGRAcDTKEJX2q07uw7OBvF
XceqrrgIEitbr0shdvCYCflQYX8HmCDxOM0ENar1ZzLE6dJm+/u9H3uOQrP7H1X7
F3JBBEgFkf6YAUsVY3eAzw7sOlwb0qIzvZinasB4c6Gx4XogFLy67hcrE9haizK6
GXgE1l5FwsLVghavMlgjnIbhZE9qZktV8RRvLOt9eHBeDyR1pdH5ap+X4HzTrxZK
eFWRz+WbcAmClo4Rs4yR1tjT8vWqyjSASy9/0xdMvjfdseCHf4cjGXt0oYIxzKL6
9S7K/ndc0EPH5HbNM58dx+vPFaqYf1oTyEeKdl+MBhJM+56luVjbdvEzdvOamCmQ
nCi6bORFmOfUHIcEU27nTnUafqXOjbME4wV/FDOKFQmzyWCCrritWgsItbLZZYtJ
BIBCu6qdgDf8kQ9Lb4/GTVNYmptpUbJ9Z9EfQgxqLcFFnoL0Iq3fuxIVQaZX6xp9
kubRLUYhv+R0pPH6LhNvWZC0LqdMiW/c08JK7WLt/sWh79JqH6j5APB09W53l8ep
ZIYQUNAeo3mQRuwB4nS0QyqodoNg0IszUAOMV+mQ87Af055k7dz18x4xOsrVWJ34
nUUHcojN5VWEoPUauU7tPkscE0O7iHGOXAM1ABYSkhXCLstkeyNEpYUEPW6v9G2V
zpDxjrJjKi5g6WckPBdwYap/xW01KfHCBRc26G28sgZCPsQdz1AVU0RrOTOWgUVu
Y5HGQUi9YUx+1RySSoSVUR6xYM8cW7YWXOp9nn/LHl0yY/O98+XTEyDufgLdJFLZ
K72fSn6zam1FH+Zg35fTcW4SSmugeJDvV7TSMxs1/oj5cV2JjUlYs7hrJY7bROtT
YSaD+QGMjcpOKykLAW0WPRwdi9cHT+IdoTJy8bc3jYAKIyWsBz2IspA9LCTQPVR2
P63kHr0iuO3NdNxxcaFVcO545nF1Ucc4upA6YEeB1gDuhricsXMfqVdFPs4UcvBs
9meXHcuqOIcns7AGeHvvZEIGm0286zRpDT229JDIq3L4y0Pe01DLgxQzfGPCtGw4
7syquw3uxfGwPuLVza2EaWFkx1eom++d4gt/llmlcgtT3/bElNWEPjNB8AZpnAQV
pyDf8OWPIMW3iX2XybC7c7XokEpQj6yNZ5ulW1cTWLDaOhh5U+2G6/ubto3kS+O/
ylTiQsgOqUVD4Xiq6bPoJQ==
`pragma protect end_protected
