// address_decode.v

// Generated using ACDS version 18.1 222

`timescale 1 ps / 1 ps
module address_decode (
		input  wire        clk_csr_clk,                                                 //                                         clk_csr.clk
		input  wire        csr_reset_n,                                                 //                                             csr.reset_n
		output wire [11:0] eth_gen_mon_0_avalon_anti_slave_0_address,                   //               eth_gen_mon_0_avalon_anti_slave_0.address
		output wire        eth_gen_mon_0_avalon_anti_slave_0_write,                     //                                                .write
		output wire        eth_gen_mon_0_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] eth_gen_mon_0_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] eth_gen_mon_0_avalon_anti_slave_0_writedata,                 //                                                .writedata
		input  wire        eth_gen_mon_0_avalon_anti_slave_0_waitrequest,               //                                                .waitrequest
		output wire [11:0] eth_gen_mon_1_avalon_anti_slave_0_address,                   //               eth_gen_mon_1_avalon_anti_slave_0.address
		output wire        eth_gen_mon_1_avalon_anti_slave_0_write,                     //                                                .write
		output wire        eth_gen_mon_1_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] eth_gen_mon_1_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] eth_gen_mon_1_avalon_anti_slave_0_writedata,                 //                                                .writedata
		input  wire        eth_gen_mon_1_avalon_anti_slave_0_waitrequest,               //                                                .waitrequest
		output wire [11:0] eth_gen_mon_10_avalon_anti_slave_0_address,                  //              eth_gen_mon_10_avalon_anti_slave_0.address
		output wire        eth_gen_mon_10_avalon_anti_slave_0_write,                    //                                                .write
		output wire        eth_gen_mon_10_avalon_anti_slave_0_read,                     //                                                .read
		input  wire [31:0] eth_gen_mon_10_avalon_anti_slave_0_readdata,                 //                                                .readdata
		output wire [31:0] eth_gen_mon_10_avalon_anti_slave_0_writedata,                //                                                .writedata
		input  wire        eth_gen_mon_10_avalon_anti_slave_0_waitrequest,              //                                                .waitrequest
		output wire [11:0] eth_gen_mon_11_avalon_anti_slave_0_address,                  //              eth_gen_mon_11_avalon_anti_slave_0.address
		output wire        eth_gen_mon_11_avalon_anti_slave_0_write,                    //                                                .write
		output wire        eth_gen_mon_11_avalon_anti_slave_0_read,                     //                                                .read
		input  wire [31:0] eth_gen_mon_11_avalon_anti_slave_0_readdata,                 //                                                .readdata
		output wire [31:0] eth_gen_mon_11_avalon_anti_slave_0_writedata,                //                                                .writedata
		input  wire        eth_gen_mon_11_avalon_anti_slave_0_waitrequest,              //                                                .waitrequest
		output wire [11:0] eth_gen_mon_2_avalon_anti_slave_0_address,                   //               eth_gen_mon_2_avalon_anti_slave_0.address
		output wire        eth_gen_mon_2_avalon_anti_slave_0_write,                     //                                                .write
		output wire        eth_gen_mon_2_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] eth_gen_mon_2_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] eth_gen_mon_2_avalon_anti_slave_0_writedata,                 //                                                .writedata
		input  wire        eth_gen_mon_2_avalon_anti_slave_0_waitrequest,               //                                                .waitrequest
		output wire [11:0] eth_gen_mon_3_avalon_anti_slave_0_address,                   //               eth_gen_mon_3_avalon_anti_slave_0.address
		output wire        eth_gen_mon_3_avalon_anti_slave_0_write,                     //                                                .write
		output wire        eth_gen_mon_3_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] eth_gen_mon_3_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] eth_gen_mon_3_avalon_anti_slave_0_writedata,                 //                                                .writedata
		input  wire        eth_gen_mon_3_avalon_anti_slave_0_waitrequest,               //                                                .waitrequest
		output wire [11:0] eth_gen_mon_4_avalon_anti_slave_0_address,                   //               eth_gen_mon_4_avalon_anti_slave_0.address
		output wire        eth_gen_mon_4_avalon_anti_slave_0_write,                     //                                                .write
		output wire        eth_gen_mon_4_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] eth_gen_mon_4_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] eth_gen_mon_4_avalon_anti_slave_0_writedata,                 //                                                .writedata
		input  wire        eth_gen_mon_4_avalon_anti_slave_0_waitrequest,               //                                                .waitrequest
		output wire [11:0] eth_gen_mon_5_avalon_anti_slave_0_address,                   //               eth_gen_mon_5_avalon_anti_slave_0.address
		output wire        eth_gen_mon_5_avalon_anti_slave_0_write,                     //                                                .write
		output wire        eth_gen_mon_5_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] eth_gen_mon_5_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] eth_gen_mon_5_avalon_anti_slave_0_writedata,                 //                                                .writedata
		input  wire        eth_gen_mon_5_avalon_anti_slave_0_waitrequest,               //                                                .waitrequest
		output wire [11:0] eth_gen_mon_6_avalon_anti_slave_0_address,                   //               eth_gen_mon_6_avalon_anti_slave_0.address
		output wire        eth_gen_mon_6_avalon_anti_slave_0_write,                     //                                                .write
		output wire        eth_gen_mon_6_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] eth_gen_mon_6_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] eth_gen_mon_6_avalon_anti_slave_0_writedata,                 //                                                .writedata
		input  wire        eth_gen_mon_6_avalon_anti_slave_0_waitrequest,               //                                                .waitrequest
		output wire [11:0] eth_gen_mon_7_avalon_anti_slave_0_address,                   //               eth_gen_mon_7_avalon_anti_slave_0.address
		output wire        eth_gen_mon_7_avalon_anti_slave_0_write,                     //                                                .write
		output wire        eth_gen_mon_7_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] eth_gen_mon_7_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] eth_gen_mon_7_avalon_anti_slave_0_writedata,                 //                                                .writedata
		input  wire        eth_gen_mon_7_avalon_anti_slave_0_waitrequest,               //                                                .waitrequest
		output wire [11:0] eth_gen_mon_8_avalon_anti_slave_0_address,                   //               eth_gen_mon_8_avalon_anti_slave_0.address
		output wire        eth_gen_mon_8_avalon_anti_slave_0_write,                     //                                                .write
		output wire        eth_gen_mon_8_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] eth_gen_mon_8_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] eth_gen_mon_8_avalon_anti_slave_0_writedata,                 //                                                .writedata
		input  wire        eth_gen_mon_8_avalon_anti_slave_0_waitrequest,               //                                                .waitrequest
		output wire [11:0] eth_gen_mon_9_avalon_anti_slave_0_address,                   //               eth_gen_mon_9_avalon_anti_slave_0.address
		output wire        eth_gen_mon_9_avalon_anti_slave_0_write,                     //                                                .write
		output wire        eth_gen_mon_9_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] eth_gen_mon_9_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] eth_gen_mon_9_avalon_anti_slave_0_writedata,                 //                                                .writedata
		input  wire        eth_gen_mon_9_avalon_anti_slave_0_waitrequest,               //                                                .waitrequest
		input  wire [15:0] merlin_master_translator_0_avalon_anti_master_0_address,     // merlin_master_translator_0_avalon_anti_master_0.address
		output wire        merlin_master_translator_0_avalon_anti_master_0_waitrequest, //                                                .waitrequest
		input  wire        merlin_master_translator_0_avalon_anti_master_0_read,        //                                                .read
		output wire [31:0] merlin_master_translator_0_avalon_anti_master_0_readdata,    //                                                .readdata
		input  wire        merlin_master_translator_0_avalon_anti_master_0_write,       //                                                .write
		input  wire [31:0] merlin_master_translator_0_avalon_anti_master_0_writedata,   //                                                .writedata
		output wire [12:0] mac_0_avalon_anti_slave_0_address,                           //                       mac_0_avalon_anti_slave_0.address
		output wire        mac_0_avalon_anti_slave_0_write,                             //                                                .write
		output wire        mac_0_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] mac_0_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] mac_0_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        mac_0_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [12:0] mac_1_avalon_anti_slave_0_address,                           //                       mac_1_avalon_anti_slave_0.address
		output wire        mac_1_avalon_anti_slave_0_write,                             //                                                .write
		output wire        mac_1_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] mac_1_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] mac_1_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        mac_1_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [12:0] mac_10_avalon_anti_slave_0_address,                          //                      mac_10_avalon_anti_slave_0.address
		output wire        mac_10_avalon_anti_slave_0_write,                            //                                                .write
		output wire        mac_10_avalon_anti_slave_0_read,                             //                                                .read
		input  wire [31:0] mac_10_avalon_anti_slave_0_readdata,                         //                                                .readdata
		output wire [31:0] mac_10_avalon_anti_slave_0_writedata,                        //                                                .writedata
		input  wire        mac_10_avalon_anti_slave_0_waitrequest,                      //                                                .waitrequest
		output wire [12:0] mac_11_avalon_anti_slave_0_address,                          //                      mac_11_avalon_anti_slave_0.address
		output wire        mac_11_avalon_anti_slave_0_write,                            //                                                .write
		output wire        mac_11_avalon_anti_slave_0_read,                             //                                                .read
		input  wire [31:0] mac_11_avalon_anti_slave_0_readdata,                         //                                                .readdata
		output wire [31:0] mac_11_avalon_anti_slave_0_writedata,                        //                                                .writedata
		input  wire        mac_11_avalon_anti_slave_0_waitrequest,                      //                                                .waitrequest
		output wire [12:0] mac_2_avalon_anti_slave_0_address,                           //                       mac_2_avalon_anti_slave_0.address
		output wire        mac_2_avalon_anti_slave_0_write,                             //                                                .write
		output wire        mac_2_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] mac_2_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] mac_2_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        mac_2_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [12:0] mac_3_avalon_anti_slave_0_address,                           //                       mac_3_avalon_anti_slave_0.address
		output wire        mac_3_avalon_anti_slave_0_write,                             //                                                .write
		output wire        mac_3_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] mac_3_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] mac_3_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        mac_3_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [12:0] mac_4_avalon_anti_slave_0_address,                           //                       mac_4_avalon_anti_slave_0.address
		output wire        mac_4_avalon_anti_slave_0_write,                             //                                                .write
		output wire        mac_4_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] mac_4_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] mac_4_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        mac_4_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [12:0] mac_5_avalon_anti_slave_0_address,                           //                       mac_5_avalon_anti_slave_0.address
		output wire        mac_5_avalon_anti_slave_0_write,                             //                                                .write
		output wire        mac_5_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] mac_5_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] mac_5_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        mac_5_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [12:0] mac_6_avalon_anti_slave_0_address,                           //                       mac_6_avalon_anti_slave_0.address
		output wire        mac_6_avalon_anti_slave_0_write,                             //                                                .write
		output wire        mac_6_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] mac_6_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] mac_6_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        mac_6_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [12:0] mac_7_avalon_anti_slave_0_address,                           //                       mac_7_avalon_anti_slave_0.address
		output wire        mac_7_avalon_anti_slave_0_write,                             //                                                .write
		output wire        mac_7_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] mac_7_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] mac_7_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        mac_7_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [12:0] mac_8_avalon_anti_slave_0_address,                           //                       mac_8_avalon_anti_slave_0.address
		output wire        mac_8_avalon_anti_slave_0_write,                             //                                                .write
		output wire        mac_8_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] mac_8_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] mac_8_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        mac_8_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [12:0] mac_9_avalon_anti_slave_0_address,                           //                       mac_9_avalon_anti_slave_0.address
		output wire        mac_9_avalon_anti_slave_0_write,                             //                                                .write
		output wire        mac_9_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] mac_9_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] mac_9_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        mac_9_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [10:0] phy_0_avalon_anti_slave_0_address,                           //                       phy_0_avalon_anti_slave_0.address
		output wire        phy_0_avalon_anti_slave_0_write,                             //                                                .write
		output wire        phy_0_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] phy_0_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] phy_0_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        phy_0_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [10:0] phy_1_avalon_anti_slave_0_address,                           //                       phy_1_avalon_anti_slave_0.address
		output wire        phy_1_avalon_anti_slave_0_write,                             //                                                .write
		output wire        phy_1_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] phy_1_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] phy_1_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        phy_1_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [10:0] phy_10_avalon_anti_slave_0_address,                          //                      phy_10_avalon_anti_slave_0.address
		output wire        phy_10_avalon_anti_slave_0_write,                            //                                                .write
		output wire        phy_10_avalon_anti_slave_0_read,                             //                                                .read
		input  wire [31:0] phy_10_avalon_anti_slave_0_readdata,                         //                                                .readdata
		output wire [31:0] phy_10_avalon_anti_slave_0_writedata,                        //                                                .writedata
		input  wire        phy_10_avalon_anti_slave_0_waitrequest,                      //                                                .waitrequest
		output wire [10:0] phy_11_avalon_anti_slave_0_address,                          //                      phy_11_avalon_anti_slave_0.address
		output wire        phy_11_avalon_anti_slave_0_write,                            //                                                .write
		output wire        phy_11_avalon_anti_slave_0_read,                             //                                                .read
		input  wire [31:0] phy_11_avalon_anti_slave_0_readdata,                         //                                                .readdata
		output wire [31:0] phy_11_avalon_anti_slave_0_writedata,                        //                                                .writedata
		input  wire        phy_11_avalon_anti_slave_0_waitrequest,                      //                                                .waitrequest
		output wire [10:0] phy_2_avalon_anti_slave_0_address,                           //                       phy_2_avalon_anti_slave_0.address
		output wire        phy_2_avalon_anti_slave_0_write,                             //                                                .write
		output wire        phy_2_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] phy_2_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] phy_2_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        phy_2_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [10:0] phy_3_avalon_anti_slave_0_address,                           //                       phy_3_avalon_anti_slave_0.address
		output wire        phy_3_avalon_anti_slave_0_write,                             //                                                .write
		output wire        phy_3_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] phy_3_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] phy_3_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        phy_3_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [10:0] phy_4_avalon_anti_slave_0_address,                           //                       phy_4_avalon_anti_slave_0.address
		output wire        phy_4_avalon_anti_slave_0_write,                             //                                                .write
		output wire        phy_4_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] phy_4_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] phy_4_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        phy_4_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [10:0] phy_5_avalon_anti_slave_0_address,                           //                       phy_5_avalon_anti_slave_0.address
		output wire        phy_5_avalon_anti_slave_0_write,                             //                                                .write
		output wire        phy_5_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] phy_5_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] phy_5_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        phy_5_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [10:0] phy_6_avalon_anti_slave_0_address,                           //                       phy_6_avalon_anti_slave_0.address
		output wire        phy_6_avalon_anti_slave_0_write,                             //                                                .write
		output wire        phy_6_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] phy_6_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] phy_6_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        phy_6_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [10:0] phy_7_avalon_anti_slave_0_address,                           //                       phy_7_avalon_anti_slave_0.address
		output wire        phy_7_avalon_anti_slave_0_write,                             //                                                .write
		output wire        phy_7_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] phy_7_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] phy_7_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        phy_7_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [10:0] phy_8_avalon_anti_slave_0_address,                           //                       phy_8_avalon_anti_slave_0.address
		output wire        phy_8_avalon_anti_slave_0_write,                             //                                                .write
		output wire        phy_8_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] phy_8_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] phy_8_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        phy_8_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [10:0] phy_9_avalon_anti_slave_0_address,                           //                       phy_9_avalon_anti_slave_0.address
		output wire        phy_9_avalon_anti_slave_0_write,                             //                                                .write
		output wire        phy_9_avalon_anti_slave_0_read,                              //                                                .read
		input  wire [31:0] phy_9_avalon_anti_slave_0_readdata,                          //                                                .readdata
		output wire [31:0] phy_9_avalon_anti_slave_0_writedata,                         //                                                .writedata
		input  wire        phy_9_avalon_anti_slave_0_waitrequest,                       //                                                .waitrequest
		output wire [2:0]  rx_sc_fifo_0_avalon_anti_slave_0_address,                    //                rx_sc_fifo_0_avalon_anti_slave_0.address
		output wire        rx_sc_fifo_0_avalon_anti_slave_0_write,                      //                                                .write
		output wire        rx_sc_fifo_0_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] rx_sc_fifo_0_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] rx_sc_fifo_0_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  rx_sc_fifo_1_avalon_anti_slave_0_address,                    //                rx_sc_fifo_1_avalon_anti_slave_0.address
		output wire        rx_sc_fifo_1_avalon_anti_slave_0_write,                      //                                                .write
		output wire        rx_sc_fifo_1_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] rx_sc_fifo_1_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] rx_sc_fifo_1_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  rx_sc_fifo_10_avalon_anti_slave_0_address,                   //               rx_sc_fifo_10_avalon_anti_slave_0.address
		output wire        rx_sc_fifo_10_avalon_anti_slave_0_write,                     //                                                .write
		output wire        rx_sc_fifo_10_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] rx_sc_fifo_10_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] rx_sc_fifo_10_avalon_anti_slave_0_writedata,                 //                                                .writedata
		output wire [2:0]  rx_sc_fifo_11_avalon_anti_slave_0_address,                   //               rx_sc_fifo_11_avalon_anti_slave_0.address
		output wire        rx_sc_fifo_11_avalon_anti_slave_0_write,                     //                                                .write
		output wire        rx_sc_fifo_11_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] rx_sc_fifo_11_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] rx_sc_fifo_11_avalon_anti_slave_0_writedata,                 //                                                .writedata
		output wire [2:0]  rx_sc_fifo_2_avalon_anti_slave_0_address,                    //                rx_sc_fifo_2_avalon_anti_slave_0.address
		output wire        rx_sc_fifo_2_avalon_anti_slave_0_write,                      //                                                .write
		output wire        rx_sc_fifo_2_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] rx_sc_fifo_2_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] rx_sc_fifo_2_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  rx_sc_fifo_3_avalon_anti_slave_0_address,                    //                rx_sc_fifo_3_avalon_anti_slave_0.address
		output wire        rx_sc_fifo_3_avalon_anti_slave_0_write,                      //                                                .write
		output wire        rx_sc_fifo_3_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] rx_sc_fifo_3_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] rx_sc_fifo_3_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  rx_sc_fifo_4_avalon_anti_slave_0_address,                    //                rx_sc_fifo_4_avalon_anti_slave_0.address
		output wire        rx_sc_fifo_4_avalon_anti_slave_0_write,                      //                                                .write
		output wire        rx_sc_fifo_4_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] rx_sc_fifo_4_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] rx_sc_fifo_4_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  rx_sc_fifo_5_avalon_anti_slave_0_address,                    //                rx_sc_fifo_5_avalon_anti_slave_0.address
		output wire        rx_sc_fifo_5_avalon_anti_slave_0_write,                      //                                                .write
		output wire        rx_sc_fifo_5_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] rx_sc_fifo_5_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] rx_sc_fifo_5_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  rx_sc_fifo_6_avalon_anti_slave_0_address,                    //                rx_sc_fifo_6_avalon_anti_slave_0.address
		output wire        rx_sc_fifo_6_avalon_anti_slave_0_write,                      //                                                .write
		output wire        rx_sc_fifo_6_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] rx_sc_fifo_6_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] rx_sc_fifo_6_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  rx_sc_fifo_7_avalon_anti_slave_0_address,                    //                rx_sc_fifo_7_avalon_anti_slave_0.address
		output wire        rx_sc_fifo_7_avalon_anti_slave_0_write,                      //                                                .write
		output wire        rx_sc_fifo_7_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] rx_sc_fifo_7_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] rx_sc_fifo_7_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  rx_sc_fifo_8_avalon_anti_slave_0_address,                    //                rx_sc_fifo_8_avalon_anti_slave_0.address
		output wire        rx_sc_fifo_8_avalon_anti_slave_0_write,                      //                                                .write
		output wire        rx_sc_fifo_8_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] rx_sc_fifo_8_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] rx_sc_fifo_8_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  rx_sc_fifo_9_avalon_anti_slave_0_address,                    //                rx_sc_fifo_9_avalon_anti_slave_0.address
		output wire        rx_sc_fifo_9_avalon_anti_slave_0_write,                      //                                                .write
		output wire        rx_sc_fifo_9_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] rx_sc_fifo_9_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] rx_sc_fifo_9_avalon_anti_slave_0_writedata,                  //                                                .writedata
		input  wire        rx_xcvr_clk_clk,                                             //                                     rx_xcvr_clk.clk
		input  wire        sync_rx_rst_reset_n,                                         //                                     sync_rx_rst.reset_n
		output wire [2:0]  tx_sc_fifo_0_avalon_anti_slave_0_address,                    //                tx_sc_fifo_0_avalon_anti_slave_0.address
		output wire        tx_sc_fifo_0_avalon_anti_slave_0_write,                      //                                                .write
		output wire        tx_sc_fifo_0_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] tx_sc_fifo_0_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] tx_sc_fifo_0_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  tx_sc_fifo_1_avalon_anti_slave_0_address,                    //                tx_sc_fifo_1_avalon_anti_slave_0.address
		output wire        tx_sc_fifo_1_avalon_anti_slave_0_write,                      //                                                .write
		output wire        tx_sc_fifo_1_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] tx_sc_fifo_1_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] tx_sc_fifo_1_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  tx_sc_fifo_10_avalon_anti_slave_0_address,                   //               tx_sc_fifo_10_avalon_anti_slave_0.address
		output wire        tx_sc_fifo_10_avalon_anti_slave_0_write,                     //                                                .write
		output wire        tx_sc_fifo_10_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] tx_sc_fifo_10_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] tx_sc_fifo_10_avalon_anti_slave_0_writedata,                 //                                                .writedata
		output wire [2:0]  tx_sc_fifo_11_avalon_anti_slave_0_address,                   //               tx_sc_fifo_11_avalon_anti_slave_0.address
		output wire        tx_sc_fifo_11_avalon_anti_slave_0_write,                     //                                                .write
		output wire        tx_sc_fifo_11_avalon_anti_slave_0_read,                      //                                                .read
		input  wire [31:0] tx_sc_fifo_11_avalon_anti_slave_0_readdata,                  //                                                .readdata
		output wire [31:0] tx_sc_fifo_11_avalon_anti_slave_0_writedata,                 //                                                .writedata
		output wire [2:0]  tx_sc_fifo_2_avalon_anti_slave_0_address,                    //                tx_sc_fifo_2_avalon_anti_slave_0.address
		output wire        tx_sc_fifo_2_avalon_anti_slave_0_write,                      //                                                .write
		output wire        tx_sc_fifo_2_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] tx_sc_fifo_2_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] tx_sc_fifo_2_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  tx_sc_fifo_3_avalon_anti_slave_0_address,                    //                tx_sc_fifo_3_avalon_anti_slave_0.address
		output wire        tx_sc_fifo_3_avalon_anti_slave_0_write,                      //                                                .write
		output wire        tx_sc_fifo_3_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] tx_sc_fifo_3_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] tx_sc_fifo_3_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  tx_sc_fifo_4_avalon_anti_slave_0_address,                    //                tx_sc_fifo_4_avalon_anti_slave_0.address
		output wire        tx_sc_fifo_4_avalon_anti_slave_0_write,                      //                                                .write
		output wire        tx_sc_fifo_4_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] tx_sc_fifo_4_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] tx_sc_fifo_4_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  tx_sc_fifo_5_avalon_anti_slave_0_address,                    //                tx_sc_fifo_5_avalon_anti_slave_0.address
		output wire        tx_sc_fifo_5_avalon_anti_slave_0_write,                      //                                                .write
		output wire        tx_sc_fifo_5_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] tx_sc_fifo_5_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] tx_sc_fifo_5_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  tx_sc_fifo_6_avalon_anti_slave_0_address,                    //                tx_sc_fifo_6_avalon_anti_slave_0.address
		output wire        tx_sc_fifo_6_avalon_anti_slave_0_write,                      //                                                .write
		output wire        tx_sc_fifo_6_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] tx_sc_fifo_6_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] tx_sc_fifo_6_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  tx_sc_fifo_7_avalon_anti_slave_0_address,                    //                tx_sc_fifo_7_avalon_anti_slave_0.address
		output wire        tx_sc_fifo_7_avalon_anti_slave_0_write,                      //                                                .write
		output wire        tx_sc_fifo_7_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] tx_sc_fifo_7_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] tx_sc_fifo_7_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  tx_sc_fifo_8_avalon_anti_slave_0_address,                    //                tx_sc_fifo_8_avalon_anti_slave_0.address
		output wire        tx_sc_fifo_8_avalon_anti_slave_0_write,                      //                                                .write
		output wire        tx_sc_fifo_8_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] tx_sc_fifo_8_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] tx_sc_fifo_8_avalon_anti_slave_0_writedata,                  //                                                .writedata
		output wire [2:0]  tx_sc_fifo_9_avalon_anti_slave_0_address,                    //                tx_sc_fifo_9_avalon_anti_slave_0.address
		output wire        tx_sc_fifo_9_avalon_anti_slave_0_write,                      //                                                .write
		output wire        tx_sc_fifo_9_avalon_anti_slave_0_read,                       //                                                .read
		input  wire [31:0] tx_sc_fifo_9_avalon_anti_slave_0_readdata,                   //                                                .readdata
		output wire [31:0] tx_sc_fifo_9_avalon_anti_slave_0_writedata,                  //                                                .writedata
		input  wire        tx_xcvr_clk_clk,                                             //                                     tx_xcvr_clk.clk
		input  wire        sync_tx_rst_reset_n,                                         //                                     sync_tx_rst.reset_n
		input  wire        tx_xcvr_half_clk_clk,                                        //                                tx_xcvr_half_clk.clk
		input  wire        sync_tx_half_rst_reset_n                                     //                                sync_tx_half_rst.reset_n
	);

	wire         clk_csr_clk_clk;                                                         // clk_csr:clk_out -> [master_0:clk_clk, merlin_master_translator_0:clk, mm_interconnect_0:clk_csr_clk_clk, mm_to_mac_0:clk, mm_to_mac_10:clk, mm_to_mac_11:clk, mm_to_mac_1:clk, mm_to_mac_2:clk, mm_to_mac_3:clk, mm_to_mac_4:clk, mm_to_mac_5:clk, mm_to_mac_6:clk, mm_to_mac_7:clk, mm_to_mac_8:clk, mm_to_mac_9:clk, mm_to_phy_0:clk, mm_to_phy_10:clk, mm_to_phy_11:clk, mm_to_phy_1:clk, mm_to_phy_2:clk, mm_to_phy_3:clk, mm_to_phy_4:clk, mm_to_phy_5:clk, mm_to_phy_6:clk, mm_to_phy_7:clk, mm_to_phy_8:clk, mm_to_phy_9:clk]
	wire         tx_xcvr_half_clk_clk_clk;                                                // tx_xcvr_half_clk:clk_out -> [eth_gen_mon_0:clk, eth_gen_mon_10:clk, eth_gen_mon_11:clk, eth_gen_mon_1:clk, eth_gen_mon_2:clk, eth_gen_mon_3:clk, eth_gen_mon_4:clk, eth_gen_mon_5:clk, eth_gen_mon_6:clk, eth_gen_mon_7:clk, eth_gen_mon_8:clk, eth_gen_mon_9:clk, mm_interconnect_0:tx_xcvr_half_clk_clk_clk, rst_controller:clk, rx_sc_fifo_0:clk, rx_sc_fifo_10:clk, rx_sc_fifo_11:clk, rx_sc_fifo_1:clk, rx_sc_fifo_2:clk, rx_sc_fifo_3:clk, rx_sc_fifo_4:clk, rx_sc_fifo_5:clk, rx_sc_fifo_6:clk, rx_sc_fifo_7:clk, rx_sc_fifo_8:clk, rx_sc_fifo_9:clk, tx_sc_fifo_0:clk, tx_sc_fifo_10:clk, tx_sc_fifo_11:clk, tx_sc_fifo_1:clk, tx_sc_fifo_2:clk, tx_sc_fifo_3:clk, tx_sc_fifo_4:clk, tx_sc_fifo_5:clk, tx_sc_fifo_6:clk, tx_sc_fifo_7:clk, tx_sc_fifo_8:clk, tx_sc_fifo_9:clk]
	wire         clk_csr_clk_reset_reset;                                                 // clk_csr:reset_n_out -> [master_0:clk_reset_reset, merlin_master_translator_0:reset, mm_interconnect_0:merlin_master_translator_0_reset_reset_bridge_in_reset_reset, mm_to_mac_0:reset, mm_to_mac_10:reset, mm_to_mac_11:reset, mm_to_mac_1:reset, mm_to_mac_2:reset, mm_to_mac_3:reset, mm_to_mac_4:reset, mm_to_mac_5:reset, mm_to_mac_6:reset, mm_to_mac_7:reset, mm_to_mac_8:reset, mm_to_mac_9:reset, mm_to_phy_0:reset, mm_to_phy_10:reset, mm_to_phy_11:reset, mm_to_phy_1:reset, mm_to_phy_2:reset, mm_to_phy_3:reset, mm_to_phy_4:reset, mm_to_phy_5:reset, mm_to_phy_6:reset, mm_to_phy_7:reset, mm_to_phy_8:reset, mm_to_phy_9:reset]
	wire         merlin_master_translator_0_avalon_universal_master_0_waitrequest;        // mm_interconnect_0:merlin_master_translator_0_avalon_universal_master_0_waitrequest -> merlin_master_translator_0:uav_waitrequest
	wire  [31:0] merlin_master_translator_0_avalon_universal_master_0_readdata;           // mm_interconnect_0:merlin_master_translator_0_avalon_universal_master_0_readdata -> merlin_master_translator_0:uav_readdata
	wire         merlin_master_translator_0_avalon_universal_master_0_debugaccess;        // merlin_master_translator_0:uav_debugaccess -> mm_interconnect_0:merlin_master_translator_0_avalon_universal_master_0_debugaccess
	wire  [31:0] merlin_master_translator_0_avalon_universal_master_0_address;            // merlin_master_translator_0:uav_address -> mm_interconnect_0:merlin_master_translator_0_avalon_universal_master_0_address
	wire         merlin_master_translator_0_avalon_universal_master_0_read;               // merlin_master_translator_0:uav_read -> mm_interconnect_0:merlin_master_translator_0_avalon_universal_master_0_read
	wire   [3:0] merlin_master_translator_0_avalon_universal_master_0_byteenable;         // merlin_master_translator_0:uav_byteenable -> mm_interconnect_0:merlin_master_translator_0_avalon_universal_master_0_byteenable
	wire         merlin_master_translator_0_avalon_universal_master_0_readdatavalid;      // mm_interconnect_0:merlin_master_translator_0_avalon_universal_master_0_readdatavalid -> merlin_master_translator_0:uav_readdatavalid
	wire         merlin_master_translator_0_avalon_universal_master_0_lock;               // merlin_master_translator_0:uav_lock -> mm_interconnect_0:merlin_master_translator_0_avalon_universal_master_0_lock
	wire         merlin_master_translator_0_avalon_universal_master_0_write;              // merlin_master_translator_0:uav_write -> mm_interconnect_0:merlin_master_translator_0_avalon_universal_master_0_write
	wire  [31:0] merlin_master_translator_0_avalon_universal_master_0_writedata;          // merlin_master_translator_0:uav_writedata -> mm_interconnect_0:merlin_master_translator_0_avalon_universal_master_0_writedata
	wire   [9:0] merlin_master_translator_0_avalon_universal_master_0_burstcount;         // merlin_master_translator_0:uav_burstcount -> mm_interconnect_0:merlin_master_translator_0_avalon_universal_master_0_burstcount
	wire  [31:0] master_0_master_readdata;                                                // mm_interconnect_0:master_0_master_readdata -> master_0:master_readdata
	wire         master_0_master_waitrequest;                                             // mm_interconnect_0:master_0_master_waitrequest -> master_0:master_waitrequest
	wire  [31:0] master_0_master_address;                                                 // master_0:master_address -> mm_interconnect_0:master_0_master_address
	wire         master_0_master_read;                                                    // master_0:master_read -> mm_interconnect_0:master_0_master_read
	wire   [3:0] master_0_master_byteenable;                                              // master_0:master_byteenable -> mm_interconnect_0:master_0_master_byteenable
	wire         master_0_master_readdatavalid;                                           // mm_interconnect_0:master_0_master_readdatavalid -> master_0:master_readdatavalid
	wire         master_0_master_write;                                                   // master_0:master_write -> mm_interconnect_0:master_0_master_write
	wire  [31:0] master_0_master_writedata;                                               // master_0:master_writedata -> mm_interconnect_0:master_0_master_writedata
	wire  [31:0] mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_readdata;         // mm_to_mac_0:uav_readdata -> mm_interconnect_0:mm_to_mac_0_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_waitrequest;      // mm_to_mac_0:uav_waitrequest -> mm_interconnect_0:mm_to_mac_0_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_mac_0_avalon_universal_slave_0_debugaccess -> mm_to_mac_0:uav_debugaccess
	wire  [14:0] mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_mac_0_avalon_universal_slave_0_address -> mm_to_mac_0:uav_address
	wire         mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_mac_0_avalon_universal_slave_0_read -> mm_to_mac_0:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_mac_0_avalon_universal_slave_0_byteenable -> mm_to_mac_0:uav_byteenable
	wire         mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_readdatavalid;    // mm_to_mac_0:uav_readdatavalid -> mm_interconnect_0:mm_to_mac_0_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_mac_0_avalon_universal_slave_0_lock -> mm_to_mac_0:uav_lock
	wire         mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_mac_0_avalon_universal_slave_0_write -> mm_to_mac_0:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_mac_0_avalon_universal_slave_0_writedata -> mm_to_mac_0:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_mac_0_avalon_universal_slave_0_burstcount -> mm_to_mac_0:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_readdata;         // mm_to_phy_0:uav_readdata -> mm_interconnect_0:mm_to_phy_0_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_waitrequest;      // mm_to_phy_0:uav_waitrequest -> mm_interconnect_0:mm_to_phy_0_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_phy_0_avalon_universal_slave_0_debugaccess -> mm_to_phy_0:uav_debugaccess
	wire  [12:0] mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_phy_0_avalon_universal_slave_0_address -> mm_to_phy_0:uav_address
	wire         mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_phy_0_avalon_universal_slave_0_read -> mm_to_phy_0:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_phy_0_avalon_universal_slave_0_byteenable -> mm_to_phy_0:uav_byteenable
	wire         mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_readdatavalid;    // mm_to_phy_0:uav_readdatavalid -> mm_interconnect_0:mm_to_phy_0_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_phy_0_avalon_universal_slave_0_lock -> mm_to_phy_0:uav_lock
	wire         mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_phy_0_avalon_universal_slave_0_write -> mm_to_phy_0:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_phy_0_avalon_universal_slave_0_writedata -> mm_to_phy_0:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_phy_0_avalon_universal_slave_0_burstcount -> mm_to_phy_0:uav_burstcount
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_readdata;        // tx_sc_fifo_0:uav_readdata -> mm_interconnect_0:tx_sc_fifo_0_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_waitrequest;     // tx_sc_fifo_0:uav_waitrequest -> mm_interconnect_0:tx_sc_fifo_0_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:tx_sc_fifo_0_avalon_universal_slave_0_debugaccess -> tx_sc_fifo_0:uav_debugaccess
	wire   [4:0] mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_address;         // mm_interconnect_0:tx_sc_fifo_0_avalon_universal_slave_0_address -> tx_sc_fifo_0:uav_address
	wire         mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_read;            // mm_interconnect_0:tx_sc_fifo_0_avalon_universal_slave_0_read -> tx_sc_fifo_0:uav_read
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:tx_sc_fifo_0_avalon_universal_slave_0_byteenable -> tx_sc_fifo_0:uav_byteenable
	wire         mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_readdatavalid;   // tx_sc_fifo_0:uav_readdatavalid -> mm_interconnect_0:tx_sc_fifo_0_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_lock;            // mm_interconnect_0:tx_sc_fifo_0_avalon_universal_slave_0_lock -> tx_sc_fifo_0:uav_lock
	wire         mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_write;           // mm_interconnect_0:tx_sc_fifo_0_avalon_universal_slave_0_write -> tx_sc_fifo_0:uav_write
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_writedata;       // mm_interconnect_0:tx_sc_fifo_0_avalon_universal_slave_0_writedata -> tx_sc_fifo_0:uav_writedata
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:tx_sc_fifo_0_avalon_universal_slave_0_burstcount -> tx_sc_fifo_0:uav_burstcount
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_readdata;        // rx_sc_fifo_0:uav_readdata -> mm_interconnect_0:rx_sc_fifo_0_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_waitrequest;     // rx_sc_fifo_0:uav_waitrequest -> mm_interconnect_0:rx_sc_fifo_0_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:rx_sc_fifo_0_avalon_universal_slave_0_debugaccess -> rx_sc_fifo_0:uav_debugaccess
	wire   [4:0] mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_address;         // mm_interconnect_0:rx_sc_fifo_0_avalon_universal_slave_0_address -> rx_sc_fifo_0:uav_address
	wire         mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_read;            // mm_interconnect_0:rx_sc_fifo_0_avalon_universal_slave_0_read -> rx_sc_fifo_0:uav_read
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:rx_sc_fifo_0_avalon_universal_slave_0_byteenable -> rx_sc_fifo_0:uav_byteenable
	wire         mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_readdatavalid;   // rx_sc_fifo_0:uav_readdatavalid -> mm_interconnect_0:rx_sc_fifo_0_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_lock;            // mm_interconnect_0:rx_sc_fifo_0_avalon_universal_slave_0_lock -> rx_sc_fifo_0:uav_lock
	wire         mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_write;           // mm_interconnect_0:rx_sc_fifo_0_avalon_universal_slave_0_write -> rx_sc_fifo_0:uav_write
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_writedata;       // mm_interconnect_0:rx_sc_fifo_0_avalon_universal_slave_0_writedata -> rx_sc_fifo_0:uav_writedata
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:rx_sc_fifo_0_avalon_universal_slave_0_burstcount -> rx_sc_fifo_0:uav_burstcount
	wire  [31:0] mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_readdata;       // eth_gen_mon_0:uav_readdata -> mm_interconnect_0:eth_gen_mon_0_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_waitrequest;    // eth_gen_mon_0:uav_waitrequest -> mm_interconnect_0:eth_gen_mon_0_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:eth_gen_mon_0_avalon_universal_slave_0_debugaccess -> eth_gen_mon_0:uav_debugaccess
	wire  [13:0] mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_address;        // mm_interconnect_0:eth_gen_mon_0_avalon_universal_slave_0_address -> eth_gen_mon_0:uav_address
	wire         mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_read;           // mm_interconnect_0:eth_gen_mon_0_avalon_universal_slave_0_read -> eth_gen_mon_0:uav_read
	wire   [3:0] mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:eth_gen_mon_0_avalon_universal_slave_0_byteenable -> eth_gen_mon_0:uav_byteenable
	wire         mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_readdatavalid;  // eth_gen_mon_0:uav_readdatavalid -> mm_interconnect_0:eth_gen_mon_0_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_lock;           // mm_interconnect_0:eth_gen_mon_0_avalon_universal_slave_0_lock -> eth_gen_mon_0:uav_lock
	wire         mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_write;          // mm_interconnect_0:eth_gen_mon_0_avalon_universal_slave_0_write -> eth_gen_mon_0:uav_write
	wire  [31:0] mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_writedata;      // mm_interconnect_0:eth_gen_mon_0_avalon_universal_slave_0_writedata -> eth_gen_mon_0:uav_writedata
	wire   [3:0] mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:eth_gen_mon_0_avalon_universal_slave_0_burstcount -> eth_gen_mon_0:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_readdata;         // mm_to_mac_1:uav_readdata -> mm_interconnect_0:mm_to_mac_1_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_waitrequest;      // mm_to_mac_1:uav_waitrequest -> mm_interconnect_0:mm_to_mac_1_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_mac_1_avalon_universal_slave_0_debugaccess -> mm_to_mac_1:uav_debugaccess
	wire  [14:0] mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_mac_1_avalon_universal_slave_0_address -> mm_to_mac_1:uav_address
	wire         mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_mac_1_avalon_universal_slave_0_read -> mm_to_mac_1:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_mac_1_avalon_universal_slave_0_byteenable -> mm_to_mac_1:uav_byteenable
	wire         mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_readdatavalid;    // mm_to_mac_1:uav_readdatavalid -> mm_interconnect_0:mm_to_mac_1_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_mac_1_avalon_universal_slave_0_lock -> mm_to_mac_1:uav_lock
	wire         mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_mac_1_avalon_universal_slave_0_write -> mm_to_mac_1:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_mac_1_avalon_universal_slave_0_writedata -> mm_to_mac_1:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_mac_1_avalon_universal_slave_0_burstcount -> mm_to_mac_1:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_readdata;         // mm_to_phy_1:uav_readdata -> mm_interconnect_0:mm_to_phy_1_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_waitrequest;      // mm_to_phy_1:uav_waitrequest -> mm_interconnect_0:mm_to_phy_1_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_phy_1_avalon_universal_slave_0_debugaccess -> mm_to_phy_1:uav_debugaccess
	wire  [12:0] mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_phy_1_avalon_universal_slave_0_address -> mm_to_phy_1:uav_address
	wire         mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_phy_1_avalon_universal_slave_0_read -> mm_to_phy_1:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_phy_1_avalon_universal_slave_0_byteenable -> mm_to_phy_1:uav_byteenable
	wire         mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_readdatavalid;    // mm_to_phy_1:uav_readdatavalid -> mm_interconnect_0:mm_to_phy_1_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_phy_1_avalon_universal_slave_0_lock -> mm_to_phy_1:uav_lock
	wire         mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_phy_1_avalon_universal_slave_0_write -> mm_to_phy_1:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_phy_1_avalon_universal_slave_0_writedata -> mm_to_phy_1:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_phy_1_avalon_universal_slave_0_burstcount -> mm_to_phy_1:uav_burstcount
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_readdata;        // rx_sc_fifo_1:uav_readdata -> mm_interconnect_0:rx_sc_fifo_1_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_waitrequest;     // rx_sc_fifo_1:uav_waitrequest -> mm_interconnect_0:rx_sc_fifo_1_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:rx_sc_fifo_1_avalon_universal_slave_0_debugaccess -> rx_sc_fifo_1:uav_debugaccess
	wire   [4:0] mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_address;         // mm_interconnect_0:rx_sc_fifo_1_avalon_universal_slave_0_address -> rx_sc_fifo_1:uav_address
	wire         mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_read;            // mm_interconnect_0:rx_sc_fifo_1_avalon_universal_slave_0_read -> rx_sc_fifo_1:uav_read
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:rx_sc_fifo_1_avalon_universal_slave_0_byteenable -> rx_sc_fifo_1:uav_byteenable
	wire         mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_readdatavalid;   // rx_sc_fifo_1:uav_readdatavalid -> mm_interconnect_0:rx_sc_fifo_1_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_lock;            // mm_interconnect_0:rx_sc_fifo_1_avalon_universal_slave_0_lock -> rx_sc_fifo_1:uav_lock
	wire         mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_write;           // mm_interconnect_0:rx_sc_fifo_1_avalon_universal_slave_0_write -> rx_sc_fifo_1:uav_write
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_writedata;       // mm_interconnect_0:rx_sc_fifo_1_avalon_universal_slave_0_writedata -> rx_sc_fifo_1:uav_writedata
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:rx_sc_fifo_1_avalon_universal_slave_0_burstcount -> rx_sc_fifo_1:uav_burstcount
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_readdata;        // tx_sc_fifo_1:uav_readdata -> mm_interconnect_0:tx_sc_fifo_1_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_waitrequest;     // tx_sc_fifo_1:uav_waitrequest -> mm_interconnect_0:tx_sc_fifo_1_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:tx_sc_fifo_1_avalon_universal_slave_0_debugaccess -> tx_sc_fifo_1:uav_debugaccess
	wire   [4:0] mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_address;         // mm_interconnect_0:tx_sc_fifo_1_avalon_universal_slave_0_address -> tx_sc_fifo_1:uav_address
	wire         mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_read;            // mm_interconnect_0:tx_sc_fifo_1_avalon_universal_slave_0_read -> tx_sc_fifo_1:uav_read
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:tx_sc_fifo_1_avalon_universal_slave_0_byteenable -> tx_sc_fifo_1:uav_byteenable
	wire         mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_readdatavalid;   // tx_sc_fifo_1:uav_readdatavalid -> mm_interconnect_0:tx_sc_fifo_1_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_lock;            // mm_interconnect_0:tx_sc_fifo_1_avalon_universal_slave_0_lock -> tx_sc_fifo_1:uav_lock
	wire         mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_write;           // mm_interconnect_0:tx_sc_fifo_1_avalon_universal_slave_0_write -> tx_sc_fifo_1:uav_write
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_writedata;       // mm_interconnect_0:tx_sc_fifo_1_avalon_universal_slave_0_writedata -> tx_sc_fifo_1:uav_writedata
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:tx_sc_fifo_1_avalon_universal_slave_0_burstcount -> tx_sc_fifo_1:uav_burstcount
	wire  [31:0] mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_readdata;       // eth_gen_mon_1:uav_readdata -> mm_interconnect_0:eth_gen_mon_1_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_waitrequest;    // eth_gen_mon_1:uav_waitrequest -> mm_interconnect_0:eth_gen_mon_1_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:eth_gen_mon_1_avalon_universal_slave_0_debugaccess -> eth_gen_mon_1:uav_debugaccess
	wire  [13:0] mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_address;        // mm_interconnect_0:eth_gen_mon_1_avalon_universal_slave_0_address -> eth_gen_mon_1:uav_address
	wire         mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_read;           // mm_interconnect_0:eth_gen_mon_1_avalon_universal_slave_0_read -> eth_gen_mon_1:uav_read
	wire   [3:0] mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:eth_gen_mon_1_avalon_universal_slave_0_byteenable -> eth_gen_mon_1:uav_byteenable
	wire         mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_readdatavalid;  // eth_gen_mon_1:uav_readdatavalid -> mm_interconnect_0:eth_gen_mon_1_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_lock;           // mm_interconnect_0:eth_gen_mon_1_avalon_universal_slave_0_lock -> eth_gen_mon_1:uav_lock
	wire         mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_write;          // mm_interconnect_0:eth_gen_mon_1_avalon_universal_slave_0_write -> eth_gen_mon_1:uav_write
	wire  [31:0] mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_writedata;      // mm_interconnect_0:eth_gen_mon_1_avalon_universal_slave_0_writedata -> eth_gen_mon_1:uav_writedata
	wire   [3:0] mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:eth_gen_mon_1_avalon_universal_slave_0_burstcount -> eth_gen_mon_1:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_readdata;         // mm_to_mac_2:uav_readdata -> mm_interconnect_0:mm_to_mac_2_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_waitrequest;      // mm_to_mac_2:uav_waitrequest -> mm_interconnect_0:mm_to_mac_2_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_mac_2_avalon_universal_slave_0_debugaccess -> mm_to_mac_2:uav_debugaccess
	wire  [14:0] mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_mac_2_avalon_universal_slave_0_address -> mm_to_mac_2:uav_address
	wire         mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_mac_2_avalon_universal_slave_0_read -> mm_to_mac_2:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_mac_2_avalon_universal_slave_0_byteenable -> mm_to_mac_2:uav_byteenable
	wire         mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_readdatavalid;    // mm_to_mac_2:uav_readdatavalid -> mm_interconnect_0:mm_to_mac_2_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_mac_2_avalon_universal_slave_0_lock -> mm_to_mac_2:uav_lock
	wire         mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_mac_2_avalon_universal_slave_0_write -> mm_to_mac_2:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_mac_2_avalon_universal_slave_0_writedata -> mm_to_mac_2:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_mac_2_avalon_universal_slave_0_burstcount -> mm_to_mac_2:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_readdata;         // mm_to_phy_2:uav_readdata -> mm_interconnect_0:mm_to_phy_2_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_waitrequest;      // mm_to_phy_2:uav_waitrequest -> mm_interconnect_0:mm_to_phy_2_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_phy_2_avalon_universal_slave_0_debugaccess -> mm_to_phy_2:uav_debugaccess
	wire  [12:0] mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_phy_2_avalon_universal_slave_0_address -> mm_to_phy_2:uav_address
	wire         mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_phy_2_avalon_universal_slave_0_read -> mm_to_phy_2:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_phy_2_avalon_universal_slave_0_byteenable -> mm_to_phy_2:uav_byteenable
	wire         mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_readdatavalid;    // mm_to_phy_2:uav_readdatavalid -> mm_interconnect_0:mm_to_phy_2_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_phy_2_avalon_universal_slave_0_lock -> mm_to_phy_2:uav_lock
	wire         mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_phy_2_avalon_universal_slave_0_write -> mm_to_phy_2:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_phy_2_avalon_universal_slave_0_writedata -> mm_to_phy_2:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_phy_2_avalon_universal_slave_0_burstcount -> mm_to_phy_2:uav_burstcount
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_readdata;        // rx_sc_fifo_2:uav_readdata -> mm_interconnect_0:rx_sc_fifo_2_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_waitrequest;     // rx_sc_fifo_2:uav_waitrequest -> mm_interconnect_0:rx_sc_fifo_2_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:rx_sc_fifo_2_avalon_universal_slave_0_debugaccess -> rx_sc_fifo_2:uav_debugaccess
	wire   [4:0] mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_address;         // mm_interconnect_0:rx_sc_fifo_2_avalon_universal_slave_0_address -> rx_sc_fifo_2:uav_address
	wire         mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_read;            // mm_interconnect_0:rx_sc_fifo_2_avalon_universal_slave_0_read -> rx_sc_fifo_2:uav_read
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:rx_sc_fifo_2_avalon_universal_slave_0_byteenable -> rx_sc_fifo_2:uav_byteenable
	wire         mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_readdatavalid;   // rx_sc_fifo_2:uav_readdatavalid -> mm_interconnect_0:rx_sc_fifo_2_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_lock;            // mm_interconnect_0:rx_sc_fifo_2_avalon_universal_slave_0_lock -> rx_sc_fifo_2:uav_lock
	wire         mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_write;           // mm_interconnect_0:rx_sc_fifo_2_avalon_universal_slave_0_write -> rx_sc_fifo_2:uav_write
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_writedata;       // mm_interconnect_0:rx_sc_fifo_2_avalon_universal_slave_0_writedata -> rx_sc_fifo_2:uav_writedata
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:rx_sc_fifo_2_avalon_universal_slave_0_burstcount -> rx_sc_fifo_2:uav_burstcount
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_readdata;        // tx_sc_fifo_2:uav_readdata -> mm_interconnect_0:tx_sc_fifo_2_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_waitrequest;     // tx_sc_fifo_2:uav_waitrequest -> mm_interconnect_0:tx_sc_fifo_2_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:tx_sc_fifo_2_avalon_universal_slave_0_debugaccess -> tx_sc_fifo_2:uav_debugaccess
	wire   [4:0] mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_address;         // mm_interconnect_0:tx_sc_fifo_2_avalon_universal_slave_0_address -> tx_sc_fifo_2:uav_address
	wire         mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_read;            // mm_interconnect_0:tx_sc_fifo_2_avalon_universal_slave_0_read -> tx_sc_fifo_2:uav_read
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:tx_sc_fifo_2_avalon_universal_slave_0_byteenable -> tx_sc_fifo_2:uav_byteenable
	wire         mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_readdatavalid;   // tx_sc_fifo_2:uav_readdatavalid -> mm_interconnect_0:tx_sc_fifo_2_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_lock;            // mm_interconnect_0:tx_sc_fifo_2_avalon_universal_slave_0_lock -> tx_sc_fifo_2:uav_lock
	wire         mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_write;           // mm_interconnect_0:tx_sc_fifo_2_avalon_universal_slave_0_write -> tx_sc_fifo_2:uav_write
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_writedata;       // mm_interconnect_0:tx_sc_fifo_2_avalon_universal_slave_0_writedata -> tx_sc_fifo_2:uav_writedata
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:tx_sc_fifo_2_avalon_universal_slave_0_burstcount -> tx_sc_fifo_2:uav_burstcount
	wire  [31:0] mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_readdata;       // eth_gen_mon_2:uav_readdata -> mm_interconnect_0:eth_gen_mon_2_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_waitrequest;    // eth_gen_mon_2:uav_waitrequest -> mm_interconnect_0:eth_gen_mon_2_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:eth_gen_mon_2_avalon_universal_slave_0_debugaccess -> eth_gen_mon_2:uav_debugaccess
	wire  [13:0] mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_address;        // mm_interconnect_0:eth_gen_mon_2_avalon_universal_slave_0_address -> eth_gen_mon_2:uav_address
	wire         mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_read;           // mm_interconnect_0:eth_gen_mon_2_avalon_universal_slave_0_read -> eth_gen_mon_2:uav_read
	wire   [3:0] mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:eth_gen_mon_2_avalon_universal_slave_0_byteenable -> eth_gen_mon_2:uav_byteenable
	wire         mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_readdatavalid;  // eth_gen_mon_2:uav_readdatavalid -> mm_interconnect_0:eth_gen_mon_2_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_lock;           // mm_interconnect_0:eth_gen_mon_2_avalon_universal_slave_0_lock -> eth_gen_mon_2:uav_lock
	wire         mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_write;          // mm_interconnect_0:eth_gen_mon_2_avalon_universal_slave_0_write -> eth_gen_mon_2:uav_write
	wire  [31:0] mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_writedata;      // mm_interconnect_0:eth_gen_mon_2_avalon_universal_slave_0_writedata -> eth_gen_mon_2:uav_writedata
	wire   [3:0] mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:eth_gen_mon_2_avalon_universal_slave_0_burstcount -> eth_gen_mon_2:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_readdata;         // mm_to_mac_3:uav_readdata -> mm_interconnect_0:mm_to_mac_3_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_waitrequest;      // mm_to_mac_3:uav_waitrequest -> mm_interconnect_0:mm_to_mac_3_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_mac_3_avalon_universal_slave_0_debugaccess -> mm_to_mac_3:uav_debugaccess
	wire  [14:0] mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_mac_3_avalon_universal_slave_0_address -> mm_to_mac_3:uav_address
	wire         mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_mac_3_avalon_universal_slave_0_read -> mm_to_mac_3:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_mac_3_avalon_universal_slave_0_byteenable -> mm_to_mac_3:uav_byteenable
	wire         mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_readdatavalid;    // mm_to_mac_3:uav_readdatavalid -> mm_interconnect_0:mm_to_mac_3_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_mac_3_avalon_universal_slave_0_lock -> mm_to_mac_3:uav_lock
	wire         mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_mac_3_avalon_universal_slave_0_write -> mm_to_mac_3:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_mac_3_avalon_universal_slave_0_writedata -> mm_to_mac_3:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_mac_3_avalon_universal_slave_0_burstcount -> mm_to_mac_3:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_readdata;         // mm_to_phy_3:uav_readdata -> mm_interconnect_0:mm_to_phy_3_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_waitrequest;      // mm_to_phy_3:uav_waitrequest -> mm_interconnect_0:mm_to_phy_3_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_phy_3_avalon_universal_slave_0_debugaccess -> mm_to_phy_3:uav_debugaccess
	wire  [12:0] mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_phy_3_avalon_universal_slave_0_address -> mm_to_phy_3:uav_address
	wire         mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_phy_3_avalon_universal_slave_0_read -> mm_to_phy_3:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_phy_3_avalon_universal_slave_0_byteenable -> mm_to_phy_3:uav_byteenable
	wire         mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_readdatavalid;    // mm_to_phy_3:uav_readdatavalid -> mm_interconnect_0:mm_to_phy_3_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_phy_3_avalon_universal_slave_0_lock -> mm_to_phy_3:uav_lock
	wire         mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_phy_3_avalon_universal_slave_0_write -> mm_to_phy_3:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_phy_3_avalon_universal_slave_0_writedata -> mm_to_phy_3:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_phy_3_avalon_universal_slave_0_burstcount -> mm_to_phy_3:uav_burstcount
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_readdata;        // rx_sc_fifo_3:uav_readdata -> mm_interconnect_0:rx_sc_fifo_3_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_waitrequest;     // rx_sc_fifo_3:uav_waitrequest -> mm_interconnect_0:rx_sc_fifo_3_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:rx_sc_fifo_3_avalon_universal_slave_0_debugaccess -> rx_sc_fifo_3:uav_debugaccess
	wire   [4:0] mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_address;         // mm_interconnect_0:rx_sc_fifo_3_avalon_universal_slave_0_address -> rx_sc_fifo_3:uav_address
	wire         mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_read;            // mm_interconnect_0:rx_sc_fifo_3_avalon_universal_slave_0_read -> rx_sc_fifo_3:uav_read
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:rx_sc_fifo_3_avalon_universal_slave_0_byteenable -> rx_sc_fifo_3:uav_byteenable
	wire         mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_readdatavalid;   // rx_sc_fifo_3:uav_readdatavalid -> mm_interconnect_0:rx_sc_fifo_3_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_lock;            // mm_interconnect_0:rx_sc_fifo_3_avalon_universal_slave_0_lock -> rx_sc_fifo_3:uav_lock
	wire         mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_write;           // mm_interconnect_0:rx_sc_fifo_3_avalon_universal_slave_0_write -> rx_sc_fifo_3:uav_write
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_writedata;       // mm_interconnect_0:rx_sc_fifo_3_avalon_universal_slave_0_writedata -> rx_sc_fifo_3:uav_writedata
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:rx_sc_fifo_3_avalon_universal_slave_0_burstcount -> rx_sc_fifo_3:uav_burstcount
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_readdata;        // tx_sc_fifo_3:uav_readdata -> mm_interconnect_0:tx_sc_fifo_3_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_waitrequest;     // tx_sc_fifo_3:uav_waitrequest -> mm_interconnect_0:tx_sc_fifo_3_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:tx_sc_fifo_3_avalon_universal_slave_0_debugaccess -> tx_sc_fifo_3:uav_debugaccess
	wire   [4:0] mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_address;         // mm_interconnect_0:tx_sc_fifo_3_avalon_universal_slave_0_address -> tx_sc_fifo_3:uav_address
	wire         mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_read;            // mm_interconnect_0:tx_sc_fifo_3_avalon_universal_slave_0_read -> tx_sc_fifo_3:uav_read
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:tx_sc_fifo_3_avalon_universal_slave_0_byteenable -> tx_sc_fifo_3:uav_byteenable
	wire         mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_readdatavalid;   // tx_sc_fifo_3:uav_readdatavalid -> mm_interconnect_0:tx_sc_fifo_3_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_lock;            // mm_interconnect_0:tx_sc_fifo_3_avalon_universal_slave_0_lock -> tx_sc_fifo_3:uav_lock
	wire         mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_write;           // mm_interconnect_0:tx_sc_fifo_3_avalon_universal_slave_0_write -> tx_sc_fifo_3:uav_write
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_writedata;       // mm_interconnect_0:tx_sc_fifo_3_avalon_universal_slave_0_writedata -> tx_sc_fifo_3:uav_writedata
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:tx_sc_fifo_3_avalon_universal_slave_0_burstcount -> tx_sc_fifo_3:uav_burstcount
	wire  [31:0] mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_readdata;       // eth_gen_mon_3:uav_readdata -> mm_interconnect_0:eth_gen_mon_3_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_waitrequest;    // eth_gen_mon_3:uav_waitrequest -> mm_interconnect_0:eth_gen_mon_3_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:eth_gen_mon_3_avalon_universal_slave_0_debugaccess -> eth_gen_mon_3:uav_debugaccess
	wire  [13:0] mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_address;        // mm_interconnect_0:eth_gen_mon_3_avalon_universal_slave_0_address -> eth_gen_mon_3:uav_address
	wire         mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_read;           // mm_interconnect_0:eth_gen_mon_3_avalon_universal_slave_0_read -> eth_gen_mon_3:uav_read
	wire   [3:0] mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:eth_gen_mon_3_avalon_universal_slave_0_byteenable -> eth_gen_mon_3:uav_byteenable
	wire         mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_readdatavalid;  // eth_gen_mon_3:uav_readdatavalid -> mm_interconnect_0:eth_gen_mon_3_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_lock;           // mm_interconnect_0:eth_gen_mon_3_avalon_universal_slave_0_lock -> eth_gen_mon_3:uav_lock
	wire         mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_write;          // mm_interconnect_0:eth_gen_mon_3_avalon_universal_slave_0_write -> eth_gen_mon_3:uav_write
	wire  [31:0] mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_writedata;      // mm_interconnect_0:eth_gen_mon_3_avalon_universal_slave_0_writedata -> eth_gen_mon_3:uav_writedata
	wire   [3:0] mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:eth_gen_mon_3_avalon_universal_slave_0_burstcount -> eth_gen_mon_3:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_readdata;         // mm_to_mac_4:uav_readdata -> mm_interconnect_0:mm_to_mac_4_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_waitrequest;      // mm_to_mac_4:uav_waitrequest -> mm_interconnect_0:mm_to_mac_4_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_mac_4_avalon_universal_slave_0_debugaccess -> mm_to_mac_4:uav_debugaccess
	wire  [14:0] mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_mac_4_avalon_universal_slave_0_address -> mm_to_mac_4:uav_address
	wire         mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_mac_4_avalon_universal_slave_0_read -> mm_to_mac_4:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_mac_4_avalon_universal_slave_0_byteenable -> mm_to_mac_4:uav_byteenable
	wire         mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_readdatavalid;    // mm_to_mac_4:uav_readdatavalid -> mm_interconnect_0:mm_to_mac_4_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_mac_4_avalon_universal_slave_0_lock -> mm_to_mac_4:uav_lock
	wire         mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_mac_4_avalon_universal_slave_0_write -> mm_to_mac_4:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_mac_4_avalon_universal_slave_0_writedata -> mm_to_mac_4:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_mac_4_avalon_universal_slave_0_burstcount -> mm_to_mac_4:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_readdata;         // mm_to_phy_4:uav_readdata -> mm_interconnect_0:mm_to_phy_4_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_waitrequest;      // mm_to_phy_4:uav_waitrequest -> mm_interconnect_0:mm_to_phy_4_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_phy_4_avalon_universal_slave_0_debugaccess -> mm_to_phy_4:uav_debugaccess
	wire  [12:0] mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_phy_4_avalon_universal_slave_0_address -> mm_to_phy_4:uav_address
	wire         mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_phy_4_avalon_universal_slave_0_read -> mm_to_phy_4:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_phy_4_avalon_universal_slave_0_byteenable -> mm_to_phy_4:uav_byteenable
	wire         mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_readdatavalid;    // mm_to_phy_4:uav_readdatavalid -> mm_interconnect_0:mm_to_phy_4_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_phy_4_avalon_universal_slave_0_lock -> mm_to_phy_4:uav_lock
	wire         mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_phy_4_avalon_universal_slave_0_write -> mm_to_phy_4:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_phy_4_avalon_universal_slave_0_writedata -> mm_to_phy_4:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_phy_4_avalon_universal_slave_0_burstcount -> mm_to_phy_4:uav_burstcount
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_readdata;        // rx_sc_fifo_4:uav_readdata -> mm_interconnect_0:rx_sc_fifo_4_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_waitrequest;     // rx_sc_fifo_4:uav_waitrequest -> mm_interconnect_0:rx_sc_fifo_4_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:rx_sc_fifo_4_avalon_universal_slave_0_debugaccess -> rx_sc_fifo_4:uav_debugaccess
	wire   [4:0] mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_address;         // mm_interconnect_0:rx_sc_fifo_4_avalon_universal_slave_0_address -> rx_sc_fifo_4:uav_address
	wire         mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_read;            // mm_interconnect_0:rx_sc_fifo_4_avalon_universal_slave_0_read -> rx_sc_fifo_4:uav_read
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:rx_sc_fifo_4_avalon_universal_slave_0_byteenable -> rx_sc_fifo_4:uav_byteenable
	wire         mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_readdatavalid;   // rx_sc_fifo_4:uav_readdatavalid -> mm_interconnect_0:rx_sc_fifo_4_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_lock;            // mm_interconnect_0:rx_sc_fifo_4_avalon_universal_slave_0_lock -> rx_sc_fifo_4:uav_lock
	wire         mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_write;           // mm_interconnect_0:rx_sc_fifo_4_avalon_universal_slave_0_write -> rx_sc_fifo_4:uav_write
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_writedata;       // mm_interconnect_0:rx_sc_fifo_4_avalon_universal_slave_0_writedata -> rx_sc_fifo_4:uav_writedata
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:rx_sc_fifo_4_avalon_universal_slave_0_burstcount -> rx_sc_fifo_4:uav_burstcount
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_readdata;        // tx_sc_fifo_4:uav_readdata -> mm_interconnect_0:tx_sc_fifo_4_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_waitrequest;     // tx_sc_fifo_4:uav_waitrequest -> mm_interconnect_0:tx_sc_fifo_4_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:tx_sc_fifo_4_avalon_universal_slave_0_debugaccess -> tx_sc_fifo_4:uav_debugaccess
	wire   [4:0] mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_address;         // mm_interconnect_0:tx_sc_fifo_4_avalon_universal_slave_0_address -> tx_sc_fifo_4:uav_address
	wire         mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_read;            // mm_interconnect_0:tx_sc_fifo_4_avalon_universal_slave_0_read -> tx_sc_fifo_4:uav_read
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:tx_sc_fifo_4_avalon_universal_slave_0_byteenable -> tx_sc_fifo_4:uav_byteenable
	wire         mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_readdatavalid;   // tx_sc_fifo_4:uav_readdatavalid -> mm_interconnect_0:tx_sc_fifo_4_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_lock;            // mm_interconnect_0:tx_sc_fifo_4_avalon_universal_slave_0_lock -> tx_sc_fifo_4:uav_lock
	wire         mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_write;           // mm_interconnect_0:tx_sc_fifo_4_avalon_universal_slave_0_write -> tx_sc_fifo_4:uav_write
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_writedata;       // mm_interconnect_0:tx_sc_fifo_4_avalon_universal_slave_0_writedata -> tx_sc_fifo_4:uav_writedata
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:tx_sc_fifo_4_avalon_universal_slave_0_burstcount -> tx_sc_fifo_4:uav_burstcount
	wire  [31:0] mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_readdata;       // eth_gen_mon_4:uav_readdata -> mm_interconnect_0:eth_gen_mon_4_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_waitrequest;    // eth_gen_mon_4:uav_waitrequest -> mm_interconnect_0:eth_gen_mon_4_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:eth_gen_mon_4_avalon_universal_slave_0_debugaccess -> eth_gen_mon_4:uav_debugaccess
	wire  [13:0] mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_address;        // mm_interconnect_0:eth_gen_mon_4_avalon_universal_slave_0_address -> eth_gen_mon_4:uav_address
	wire         mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_read;           // mm_interconnect_0:eth_gen_mon_4_avalon_universal_slave_0_read -> eth_gen_mon_4:uav_read
	wire   [3:0] mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:eth_gen_mon_4_avalon_universal_slave_0_byteenable -> eth_gen_mon_4:uav_byteenable
	wire         mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_readdatavalid;  // eth_gen_mon_4:uav_readdatavalid -> mm_interconnect_0:eth_gen_mon_4_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_lock;           // mm_interconnect_0:eth_gen_mon_4_avalon_universal_slave_0_lock -> eth_gen_mon_4:uav_lock
	wire         mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_write;          // mm_interconnect_0:eth_gen_mon_4_avalon_universal_slave_0_write -> eth_gen_mon_4:uav_write
	wire  [31:0] mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_writedata;      // mm_interconnect_0:eth_gen_mon_4_avalon_universal_slave_0_writedata -> eth_gen_mon_4:uav_writedata
	wire   [3:0] mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:eth_gen_mon_4_avalon_universal_slave_0_burstcount -> eth_gen_mon_4:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_readdata;         // mm_to_mac_5:uav_readdata -> mm_interconnect_0:mm_to_mac_5_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_waitrequest;      // mm_to_mac_5:uav_waitrequest -> mm_interconnect_0:mm_to_mac_5_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_mac_5_avalon_universal_slave_0_debugaccess -> mm_to_mac_5:uav_debugaccess
	wire  [14:0] mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_mac_5_avalon_universal_slave_0_address -> mm_to_mac_5:uav_address
	wire         mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_mac_5_avalon_universal_slave_0_read -> mm_to_mac_5:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_mac_5_avalon_universal_slave_0_byteenable -> mm_to_mac_5:uav_byteenable
	wire         mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_readdatavalid;    // mm_to_mac_5:uav_readdatavalid -> mm_interconnect_0:mm_to_mac_5_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_mac_5_avalon_universal_slave_0_lock -> mm_to_mac_5:uav_lock
	wire         mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_mac_5_avalon_universal_slave_0_write -> mm_to_mac_5:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_mac_5_avalon_universal_slave_0_writedata -> mm_to_mac_5:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_mac_5_avalon_universal_slave_0_burstcount -> mm_to_mac_5:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_readdata;         // mm_to_phy_5:uav_readdata -> mm_interconnect_0:mm_to_phy_5_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_waitrequest;      // mm_to_phy_5:uav_waitrequest -> mm_interconnect_0:mm_to_phy_5_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_phy_5_avalon_universal_slave_0_debugaccess -> mm_to_phy_5:uav_debugaccess
	wire  [12:0] mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_phy_5_avalon_universal_slave_0_address -> mm_to_phy_5:uav_address
	wire         mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_phy_5_avalon_universal_slave_0_read -> mm_to_phy_5:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_phy_5_avalon_universal_slave_0_byteenable -> mm_to_phy_5:uav_byteenable
	wire         mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_readdatavalid;    // mm_to_phy_5:uav_readdatavalid -> mm_interconnect_0:mm_to_phy_5_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_phy_5_avalon_universal_slave_0_lock -> mm_to_phy_5:uav_lock
	wire         mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_phy_5_avalon_universal_slave_0_write -> mm_to_phy_5:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_phy_5_avalon_universal_slave_0_writedata -> mm_to_phy_5:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_phy_5_avalon_universal_slave_0_burstcount -> mm_to_phy_5:uav_burstcount
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_readdata;        // rx_sc_fifo_5:uav_readdata -> mm_interconnect_0:rx_sc_fifo_5_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_waitrequest;     // rx_sc_fifo_5:uav_waitrequest -> mm_interconnect_0:rx_sc_fifo_5_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:rx_sc_fifo_5_avalon_universal_slave_0_debugaccess -> rx_sc_fifo_5:uav_debugaccess
	wire   [4:0] mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_address;         // mm_interconnect_0:rx_sc_fifo_5_avalon_universal_slave_0_address -> rx_sc_fifo_5:uav_address
	wire         mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_read;            // mm_interconnect_0:rx_sc_fifo_5_avalon_universal_slave_0_read -> rx_sc_fifo_5:uav_read
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:rx_sc_fifo_5_avalon_universal_slave_0_byteenable -> rx_sc_fifo_5:uav_byteenable
	wire         mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_readdatavalid;   // rx_sc_fifo_5:uav_readdatavalid -> mm_interconnect_0:rx_sc_fifo_5_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_lock;            // mm_interconnect_0:rx_sc_fifo_5_avalon_universal_slave_0_lock -> rx_sc_fifo_5:uav_lock
	wire         mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_write;           // mm_interconnect_0:rx_sc_fifo_5_avalon_universal_slave_0_write -> rx_sc_fifo_5:uav_write
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_writedata;       // mm_interconnect_0:rx_sc_fifo_5_avalon_universal_slave_0_writedata -> rx_sc_fifo_5:uav_writedata
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:rx_sc_fifo_5_avalon_universal_slave_0_burstcount -> rx_sc_fifo_5:uav_burstcount
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_readdata;        // tx_sc_fifo_5:uav_readdata -> mm_interconnect_0:tx_sc_fifo_5_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_waitrequest;     // tx_sc_fifo_5:uav_waitrequest -> mm_interconnect_0:tx_sc_fifo_5_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:tx_sc_fifo_5_avalon_universal_slave_0_debugaccess -> tx_sc_fifo_5:uav_debugaccess
	wire   [4:0] mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_address;         // mm_interconnect_0:tx_sc_fifo_5_avalon_universal_slave_0_address -> tx_sc_fifo_5:uav_address
	wire         mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_read;            // mm_interconnect_0:tx_sc_fifo_5_avalon_universal_slave_0_read -> tx_sc_fifo_5:uav_read
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:tx_sc_fifo_5_avalon_universal_slave_0_byteenable -> tx_sc_fifo_5:uav_byteenable
	wire         mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_readdatavalid;   // tx_sc_fifo_5:uav_readdatavalid -> mm_interconnect_0:tx_sc_fifo_5_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_lock;            // mm_interconnect_0:tx_sc_fifo_5_avalon_universal_slave_0_lock -> tx_sc_fifo_5:uav_lock
	wire         mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_write;           // mm_interconnect_0:tx_sc_fifo_5_avalon_universal_slave_0_write -> tx_sc_fifo_5:uav_write
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_writedata;       // mm_interconnect_0:tx_sc_fifo_5_avalon_universal_slave_0_writedata -> tx_sc_fifo_5:uav_writedata
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:tx_sc_fifo_5_avalon_universal_slave_0_burstcount -> tx_sc_fifo_5:uav_burstcount
	wire  [31:0] mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_readdata;       // eth_gen_mon_5:uav_readdata -> mm_interconnect_0:eth_gen_mon_5_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_waitrequest;    // eth_gen_mon_5:uav_waitrequest -> mm_interconnect_0:eth_gen_mon_5_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:eth_gen_mon_5_avalon_universal_slave_0_debugaccess -> eth_gen_mon_5:uav_debugaccess
	wire  [13:0] mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_address;        // mm_interconnect_0:eth_gen_mon_5_avalon_universal_slave_0_address -> eth_gen_mon_5:uav_address
	wire         mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_read;           // mm_interconnect_0:eth_gen_mon_5_avalon_universal_slave_0_read -> eth_gen_mon_5:uav_read
	wire   [3:0] mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:eth_gen_mon_5_avalon_universal_slave_0_byteenable -> eth_gen_mon_5:uav_byteenable
	wire         mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_readdatavalid;  // eth_gen_mon_5:uav_readdatavalid -> mm_interconnect_0:eth_gen_mon_5_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_lock;           // mm_interconnect_0:eth_gen_mon_5_avalon_universal_slave_0_lock -> eth_gen_mon_5:uav_lock
	wire         mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_write;          // mm_interconnect_0:eth_gen_mon_5_avalon_universal_slave_0_write -> eth_gen_mon_5:uav_write
	wire  [31:0] mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_writedata;      // mm_interconnect_0:eth_gen_mon_5_avalon_universal_slave_0_writedata -> eth_gen_mon_5:uav_writedata
	wire   [3:0] mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:eth_gen_mon_5_avalon_universal_slave_0_burstcount -> eth_gen_mon_5:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_readdata;         // mm_to_mac_6:uav_readdata -> mm_interconnect_0:mm_to_mac_6_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_waitrequest;      // mm_to_mac_6:uav_waitrequest -> mm_interconnect_0:mm_to_mac_6_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_mac_6_avalon_universal_slave_0_debugaccess -> mm_to_mac_6:uav_debugaccess
	wire  [14:0] mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_mac_6_avalon_universal_slave_0_address -> mm_to_mac_6:uav_address
	wire         mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_mac_6_avalon_universal_slave_0_read -> mm_to_mac_6:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_mac_6_avalon_universal_slave_0_byteenable -> mm_to_mac_6:uav_byteenable
	wire         mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_readdatavalid;    // mm_to_mac_6:uav_readdatavalid -> mm_interconnect_0:mm_to_mac_6_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_mac_6_avalon_universal_slave_0_lock -> mm_to_mac_6:uav_lock
	wire         mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_mac_6_avalon_universal_slave_0_write -> mm_to_mac_6:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_mac_6_avalon_universal_slave_0_writedata -> mm_to_mac_6:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_mac_6_avalon_universal_slave_0_burstcount -> mm_to_mac_6:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_readdata;         // mm_to_phy_6:uav_readdata -> mm_interconnect_0:mm_to_phy_6_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_waitrequest;      // mm_to_phy_6:uav_waitrequest -> mm_interconnect_0:mm_to_phy_6_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_phy_6_avalon_universal_slave_0_debugaccess -> mm_to_phy_6:uav_debugaccess
	wire  [12:0] mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_phy_6_avalon_universal_slave_0_address -> mm_to_phy_6:uav_address
	wire         mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_phy_6_avalon_universal_slave_0_read -> mm_to_phy_6:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_phy_6_avalon_universal_slave_0_byteenable -> mm_to_phy_6:uav_byteenable
	wire         mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_readdatavalid;    // mm_to_phy_6:uav_readdatavalid -> mm_interconnect_0:mm_to_phy_6_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_phy_6_avalon_universal_slave_0_lock -> mm_to_phy_6:uav_lock
	wire         mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_phy_6_avalon_universal_slave_0_write -> mm_to_phy_6:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_phy_6_avalon_universal_slave_0_writedata -> mm_to_phy_6:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_phy_6_avalon_universal_slave_0_burstcount -> mm_to_phy_6:uav_burstcount
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_readdata;        // rx_sc_fifo_6:uav_readdata -> mm_interconnect_0:rx_sc_fifo_6_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_waitrequest;     // rx_sc_fifo_6:uav_waitrequest -> mm_interconnect_0:rx_sc_fifo_6_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:rx_sc_fifo_6_avalon_universal_slave_0_debugaccess -> rx_sc_fifo_6:uav_debugaccess
	wire   [4:0] mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_address;         // mm_interconnect_0:rx_sc_fifo_6_avalon_universal_slave_0_address -> rx_sc_fifo_6:uav_address
	wire         mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_read;            // mm_interconnect_0:rx_sc_fifo_6_avalon_universal_slave_0_read -> rx_sc_fifo_6:uav_read
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:rx_sc_fifo_6_avalon_universal_slave_0_byteenable -> rx_sc_fifo_6:uav_byteenable
	wire         mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_readdatavalid;   // rx_sc_fifo_6:uav_readdatavalid -> mm_interconnect_0:rx_sc_fifo_6_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_lock;            // mm_interconnect_0:rx_sc_fifo_6_avalon_universal_slave_0_lock -> rx_sc_fifo_6:uav_lock
	wire         mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_write;           // mm_interconnect_0:rx_sc_fifo_6_avalon_universal_slave_0_write -> rx_sc_fifo_6:uav_write
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_writedata;       // mm_interconnect_0:rx_sc_fifo_6_avalon_universal_slave_0_writedata -> rx_sc_fifo_6:uav_writedata
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:rx_sc_fifo_6_avalon_universal_slave_0_burstcount -> rx_sc_fifo_6:uav_burstcount
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_readdata;        // tx_sc_fifo_6:uav_readdata -> mm_interconnect_0:tx_sc_fifo_6_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_waitrequest;     // tx_sc_fifo_6:uav_waitrequest -> mm_interconnect_0:tx_sc_fifo_6_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:tx_sc_fifo_6_avalon_universal_slave_0_debugaccess -> tx_sc_fifo_6:uav_debugaccess
	wire   [4:0] mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_address;         // mm_interconnect_0:tx_sc_fifo_6_avalon_universal_slave_0_address -> tx_sc_fifo_6:uav_address
	wire         mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_read;            // mm_interconnect_0:tx_sc_fifo_6_avalon_universal_slave_0_read -> tx_sc_fifo_6:uav_read
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:tx_sc_fifo_6_avalon_universal_slave_0_byteenable -> tx_sc_fifo_6:uav_byteenable
	wire         mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_readdatavalid;   // tx_sc_fifo_6:uav_readdatavalid -> mm_interconnect_0:tx_sc_fifo_6_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_lock;            // mm_interconnect_0:tx_sc_fifo_6_avalon_universal_slave_0_lock -> tx_sc_fifo_6:uav_lock
	wire         mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_write;           // mm_interconnect_0:tx_sc_fifo_6_avalon_universal_slave_0_write -> tx_sc_fifo_6:uav_write
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_writedata;       // mm_interconnect_0:tx_sc_fifo_6_avalon_universal_slave_0_writedata -> tx_sc_fifo_6:uav_writedata
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:tx_sc_fifo_6_avalon_universal_slave_0_burstcount -> tx_sc_fifo_6:uav_burstcount
	wire  [31:0] mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_readdata;       // eth_gen_mon_6:uav_readdata -> mm_interconnect_0:eth_gen_mon_6_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_waitrequest;    // eth_gen_mon_6:uav_waitrequest -> mm_interconnect_0:eth_gen_mon_6_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:eth_gen_mon_6_avalon_universal_slave_0_debugaccess -> eth_gen_mon_6:uav_debugaccess
	wire  [13:0] mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_address;        // mm_interconnect_0:eth_gen_mon_6_avalon_universal_slave_0_address -> eth_gen_mon_6:uav_address
	wire         mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_read;           // mm_interconnect_0:eth_gen_mon_6_avalon_universal_slave_0_read -> eth_gen_mon_6:uav_read
	wire   [3:0] mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:eth_gen_mon_6_avalon_universal_slave_0_byteenable -> eth_gen_mon_6:uav_byteenable
	wire         mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_readdatavalid;  // eth_gen_mon_6:uav_readdatavalid -> mm_interconnect_0:eth_gen_mon_6_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_lock;           // mm_interconnect_0:eth_gen_mon_6_avalon_universal_slave_0_lock -> eth_gen_mon_6:uav_lock
	wire         mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_write;          // mm_interconnect_0:eth_gen_mon_6_avalon_universal_slave_0_write -> eth_gen_mon_6:uav_write
	wire  [31:0] mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_writedata;      // mm_interconnect_0:eth_gen_mon_6_avalon_universal_slave_0_writedata -> eth_gen_mon_6:uav_writedata
	wire   [3:0] mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:eth_gen_mon_6_avalon_universal_slave_0_burstcount -> eth_gen_mon_6:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_readdata;         // mm_to_mac_7:uav_readdata -> mm_interconnect_0:mm_to_mac_7_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_waitrequest;      // mm_to_mac_7:uav_waitrequest -> mm_interconnect_0:mm_to_mac_7_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_mac_7_avalon_universal_slave_0_debugaccess -> mm_to_mac_7:uav_debugaccess
	wire  [14:0] mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_mac_7_avalon_universal_slave_0_address -> mm_to_mac_7:uav_address
	wire         mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_mac_7_avalon_universal_slave_0_read -> mm_to_mac_7:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_mac_7_avalon_universal_slave_0_byteenable -> mm_to_mac_7:uav_byteenable
	wire         mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_readdatavalid;    // mm_to_mac_7:uav_readdatavalid -> mm_interconnect_0:mm_to_mac_7_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_mac_7_avalon_universal_slave_0_lock -> mm_to_mac_7:uav_lock
	wire         mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_mac_7_avalon_universal_slave_0_write -> mm_to_mac_7:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_mac_7_avalon_universal_slave_0_writedata -> mm_to_mac_7:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_mac_7_avalon_universal_slave_0_burstcount -> mm_to_mac_7:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_readdata;         // mm_to_phy_7:uav_readdata -> mm_interconnect_0:mm_to_phy_7_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_waitrequest;      // mm_to_phy_7:uav_waitrequest -> mm_interconnect_0:mm_to_phy_7_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_phy_7_avalon_universal_slave_0_debugaccess -> mm_to_phy_7:uav_debugaccess
	wire  [12:0] mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_phy_7_avalon_universal_slave_0_address -> mm_to_phy_7:uav_address
	wire         mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_phy_7_avalon_universal_slave_0_read -> mm_to_phy_7:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_phy_7_avalon_universal_slave_0_byteenable -> mm_to_phy_7:uav_byteenable
	wire         mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_readdatavalid;    // mm_to_phy_7:uav_readdatavalid -> mm_interconnect_0:mm_to_phy_7_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_phy_7_avalon_universal_slave_0_lock -> mm_to_phy_7:uav_lock
	wire         mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_phy_7_avalon_universal_slave_0_write -> mm_to_phy_7:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_phy_7_avalon_universal_slave_0_writedata -> mm_to_phy_7:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_phy_7_avalon_universal_slave_0_burstcount -> mm_to_phy_7:uav_burstcount
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_readdata;        // rx_sc_fifo_7:uav_readdata -> mm_interconnect_0:rx_sc_fifo_7_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_waitrequest;     // rx_sc_fifo_7:uav_waitrequest -> mm_interconnect_0:rx_sc_fifo_7_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:rx_sc_fifo_7_avalon_universal_slave_0_debugaccess -> rx_sc_fifo_7:uav_debugaccess
	wire   [4:0] mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_address;         // mm_interconnect_0:rx_sc_fifo_7_avalon_universal_slave_0_address -> rx_sc_fifo_7:uav_address
	wire         mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_read;            // mm_interconnect_0:rx_sc_fifo_7_avalon_universal_slave_0_read -> rx_sc_fifo_7:uav_read
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:rx_sc_fifo_7_avalon_universal_slave_0_byteenable -> rx_sc_fifo_7:uav_byteenable
	wire         mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_readdatavalid;   // rx_sc_fifo_7:uav_readdatavalid -> mm_interconnect_0:rx_sc_fifo_7_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_lock;            // mm_interconnect_0:rx_sc_fifo_7_avalon_universal_slave_0_lock -> rx_sc_fifo_7:uav_lock
	wire         mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_write;           // mm_interconnect_0:rx_sc_fifo_7_avalon_universal_slave_0_write -> rx_sc_fifo_7:uav_write
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_writedata;       // mm_interconnect_0:rx_sc_fifo_7_avalon_universal_slave_0_writedata -> rx_sc_fifo_7:uav_writedata
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:rx_sc_fifo_7_avalon_universal_slave_0_burstcount -> rx_sc_fifo_7:uav_burstcount
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_readdata;        // tx_sc_fifo_7:uav_readdata -> mm_interconnect_0:tx_sc_fifo_7_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_waitrequest;     // tx_sc_fifo_7:uav_waitrequest -> mm_interconnect_0:tx_sc_fifo_7_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:tx_sc_fifo_7_avalon_universal_slave_0_debugaccess -> tx_sc_fifo_7:uav_debugaccess
	wire   [4:0] mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_address;         // mm_interconnect_0:tx_sc_fifo_7_avalon_universal_slave_0_address -> tx_sc_fifo_7:uav_address
	wire         mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_read;            // mm_interconnect_0:tx_sc_fifo_7_avalon_universal_slave_0_read -> tx_sc_fifo_7:uav_read
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:tx_sc_fifo_7_avalon_universal_slave_0_byteenable -> tx_sc_fifo_7:uav_byteenable
	wire         mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_readdatavalid;   // tx_sc_fifo_7:uav_readdatavalid -> mm_interconnect_0:tx_sc_fifo_7_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_lock;            // mm_interconnect_0:tx_sc_fifo_7_avalon_universal_slave_0_lock -> tx_sc_fifo_7:uav_lock
	wire         mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_write;           // mm_interconnect_0:tx_sc_fifo_7_avalon_universal_slave_0_write -> tx_sc_fifo_7:uav_write
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_writedata;       // mm_interconnect_0:tx_sc_fifo_7_avalon_universal_slave_0_writedata -> tx_sc_fifo_7:uav_writedata
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:tx_sc_fifo_7_avalon_universal_slave_0_burstcount -> tx_sc_fifo_7:uav_burstcount
	wire  [31:0] mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_readdata;       // eth_gen_mon_7:uav_readdata -> mm_interconnect_0:eth_gen_mon_7_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_waitrequest;    // eth_gen_mon_7:uav_waitrequest -> mm_interconnect_0:eth_gen_mon_7_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:eth_gen_mon_7_avalon_universal_slave_0_debugaccess -> eth_gen_mon_7:uav_debugaccess
	wire  [13:0] mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_address;        // mm_interconnect_0:eth_gen_mon_7_avalon_universal_slave_0_address -> eth_gen_mon_7:uav_address
	wire         mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_read;           // mm_interconnect_0:eth_gen_mon_7_avalon_universal_slave_0_read -> eth_gen_mon_7:uav_read
	wire   [3:0] mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:eth_gen_mon_7_avalon_universal_slave_0_byteenable -> eth_gen_mon_7:uav_byteenable
	wire         mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_readdatavalid;  // eth_gen_mon_7:uav_readdatavalid -> mm_interconnect_0:eth_gen_mon_7_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_lock;           // mm_interconnect_0:eth_gen_mon_7_avalon_universal_slave_0_lock -> eth_gen_mon_7:uav_lock
	wire         mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_write;          // mm_interconnect_0:eth_gen_mon_7_avalon_universal_slave_0_write -> eth_gen_mon_7:uav_write
	wire  [31:0] mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_writedata;      // mm_interconnect_0:eth_gen_mon_7_avalon_universal_slave_0_writedata -> eth_gen_mon_7:uav_writedata
	wire   [3:0] mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:eth_gen_mon_7_avalon_universal_slave_0_burstcount -> eth_gen_mon_7:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_readdata;         // mm_to_mac_8:uav_readdata -> mm_interconnect_0:mm_to_mac_8_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_waitrequest;      // mm_to_mac_8:uav_waitrequest -> mm_interconnect_0:mm_to_mac_8_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_mac_8_avalon_universal_slave_0_debugaccess -> mm_to_mac_8:uav_debugaccess
	wire  [14:0] mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_mac_8_avalon_universal_slave_0_address -> mm_to_mac_8:uav_address
	wire         mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_mac_8_avalon_universal_slave_0_read -> mm_to_mac_8:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_mac_8_avalon_universal_slave_0_byteenable -> mm_to_mac_8:uav_byteenable
	wire         mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_readdatavalid;    // mm_to_mac_8:uav_readdatavalid -> mm_interconnect_0:mm_to_mac_8_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_mac_8_avalon_universal_slave_0_lock -> mm_to_mac_8:uav_lock
	wire         mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_mac_8_avalon_universal_slave_0_write -> mm_to_mac_8:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_mac_8_avalon_universal_slave_0_writedata -> mm_to_mac_8:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_mac_8_avalon_universal_slave_0_burstcount -> mm_to_mac_8:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_readdata;         // mm_to_phy_8:uav_readdata -> mm_interconnect_0:mm_to_phy_8_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_waitrequest;      // mm_to_phy_8:uav_waitrequest -> mm_interconnect_0:mm_to_phy_8_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_phy_8_avalon_universal_slave_0_debugaccess -> mm_to_phy_8:uav_debugaccess
	wire  [12:0] mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_phy_8_avalon_universal_slave_0_address -> mm_to_phy_8:uav_address
	wire         mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_phy_8_avalon_universal_slave_0_read -> mm_to_phy_8:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_phy_8_avalon_universal_slave_0_byteenable -> mm_to_phy_8:uav_byteenable
	wire         mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_readdatavalid;    // mm_to_phy_8:uav_readdatavalid -> mm_interconnect_0:mm_to_phy_8_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_phy_8_avalon_universal_slave_0_lock -> mm_to_phy_8:uav_lock
	wire         mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_phy_8_avalon_universal_slave_0_write -> mm_to_phy_8:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_phy_8_avalon_universal_slave_0_writedata -> mm_to_phy_8:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_phy_8_avalon_universal_slave_0_burstcount -> mm_to_phy_8:uav_burstcount
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_readdata;        // rx_sc_fifo_8:uav_readdata -> mm_interconnect_0:rx_sc_fifo_8_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_waitrequest;     // rx_sc_fifo_8:uav_waitrequest -> mm_interconnect_0:rx_sc_fifo_8_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:rx_sc_fifo_8_avalon_universal_slave_0_debugaccess -> rx_sc_fifo_8:uav_debugaccess
	wire   [4:0] mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_address;         // mm_interconnect_0:rx_sc_fifo_8_avalon_universal_slave_0_address -> rx_sc_fifo_8:uav_address
	wire         mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_read;            // mm_interconnect_0:rx_sc_fifo_8_avalon_universal_slave_0_read -> rx_sc_fifo_8:uav_read
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:rx_sc_fifo_8_avalon_universal_slave_0_byteenable -> rx_sc_fifo_8:uav_byteenable
	wire         mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_readdatavalid;   // rx_sc_fifo_8:uav_readdatavalid -> mm_interconnect_0:rx_sc_fifo_8_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_lock;            // mm_interconnect_0:rx_sc_fifo_8_avalon_universal_slave_0_lock -> rx_sc_fifo_8:uav_lock
	wire         mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_write;           // mm_interconnect_0:rx_sc_fifo_8_avalon_universal_slave_0_write -> rx_sc_fifo_8:uav_write
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_writedata;       // mm_interconnect_0:rx_sc_fifo_8_avalon_universal_slave_0_writedata -> rx_sc_fifo_8:uav_writedata
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:rx_sc_fifo_8_avalon_universal_slave_0_burstcount -> rx_sc_fifo_8:uav_burstcount
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_readdata;        // tx_sc_fifo_8:uav_readdata -> mm_interconnect_0:tx_sc_fifo_8_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_waitrequest;     // tx_sc_fifo_8:uav_waitrequest -> mm_interconnect_0:tx_sc_fifo_8_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:tx_sc_fifo_8_avalon_universal_slave_0_debugaccess -> tx_sc_fifo_8:uav_debugaccess
	wire   [4:0] mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_address;         // mm_interconnect_0:tx_sc_fifo_8_avalon_universal_slave_0_address -> tx_sc_fifo_8:uav_address
	wire         mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_read;            // mm_interconnect_0:tx_sc_fifo_8_avalon_universal_slave_0_read -> tx_sc_fifo_8:uav_read
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:tx_sc_fifo_8_avalon_universal_slave_0_byteenable -> tx_sc_fifo_8:uav_byteenable
	wire         mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_readdatavalid;   // tx_sc_fifo_8:uav_readdatavalid -> mm_interconnect_0:tx_sc_fifo_8_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_lock;            // mm_interconnect_0:tx_sc_fifo_8_avalon_universal_slave_0_lock -> tx_sc_fifo_8:uav_lock
	wire         mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_write;           // mm_interconnect_0:tx_sc_fifo_8_avalon_universal_slave_0_write -> tx_sc_fifo_8:uav_write
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_writedata;       // mm_interconnect_0:tx_sc_fifo_8_avalon_universal_slave_0_writedata -> tx_sc_fifo_8:uav_writedata
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:tx_sc_fifo_8_avalon_universal_slave_0_burstcount -> tx_sc_fifo_8:uav_burstcount
	wire  [31:0] mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_readdata;       // eth_gen_mon_8:uav_readdata -> mm_interconnect_0:eth_gen_mon_8_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_waitrequest;    // eth_gen_mon_8:uav_waitrequest -> mm_interconnect_0:eth_gen_mon_8_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:eth_gen_mon_8_avalon_universal_slave_0_debugaccess -> eth_gen_mon_8:uav_debugaccess
	wire  [13:0] mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_address;        // mm_interconnect_0:eth_gen_mon_8_avalon_universal_slave_0_address -> eth_gen_mon_8:uav_address
	wire         mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_read;           // mm_interconnect_0:eth_gen_mon_8_avalon_universal_slave_0_read -> eth_gen_mon_8:uav_read
	wire   [3:0] mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:eth_gen_mon_8_avalon_universal_slave_0_byteenable -> eth_gen_mon_8:uav_byteenable
	wire         mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_readdatavalid;  // eth_gen_mon_8:uav_readdatavalid -> mm_interconnect_0:eth_gen_mon_8_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_lock;           // mm_interconnect_0:eth_gen_mon_8_avalon_universal_slave_0_lock -> eth_gen_mon_8:uav_lock
	wire         mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_write;          // mm_interconnect_0:eth_gen_mon_8_avalon_universal_slave_0_write -> eth_gen_mon_8:uav_write
	wire  [31:0] mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_writedata;      // mm_interconnect_0:eth_gen_mon_8_avalon_universal_slave_0_writedata -> eth_gen_mon_8:uav_writedata
	wire   [3:0] mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:eth_gen_mon_8_avalon_universal_slave_0_burstcount -> eth_gen_mon_8:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_readdata;         // mm_to_mac_9:uav_readdata -> mm_interconnect_0:mm_to_mac_9_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_waitrequest;      // mm_to_mac_9:uav_waitrequest -> mm_interconnect_0:mm_to_mac_9_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_mac_9_avalon_universal_slave_0_debugaccess -> mm_to_mac_9:uav_debugaccess
	wire  [14:0] mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_mac_9_avalon_universal_slave_0_address -> mm_to_mac_9:uav_address
	wire         mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_mac_9_avalon_universal_slave_0_read -> mm_to_mac_9:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_mac_9_avalon_universal_slave_0_byteenable -> mm_to_mac_9:uav_byteenable
	wire         mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_readdatavalid;    // mm_to_mac_9:uav_readdatavalid -> mm_interconnect_0:mm_to_mac_9_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_mac_9_avalon_universal_slave_0_lock -> mm_to_mac_9:uav_lock
	wire         mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_mac_9_avalon_universal_slave_0_write -> mm_to_mac_9:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_mac_9_avalon_universal_slave_0_writedata -> mm_to_mac_9:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_mac_9_avalon_universal_slave_0_burstcount -> mm_to_mac_9:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_readdata;         // mm_to_phy_9:uav_readdata -> mm_interconnect_0:mm_to_phy_9_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_waitrequest;      // mm_to_phy_9:uav_waitrequest -> mm_interconnect_0:mm_to_phy_9_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_debugaccess;      // mm_interconnect_0:mm_to_phy_9_avalon_universal_slave_0_debugaccess -> mm_to_phy_9:uav_debugaccess
	wire  [12:0] mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_address;          // mm_interconnect_0:mm_to_phy_9_avalon_universal_slave_0_address -> mm_to_phy_9:uav_address
	wire         mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_read;             // mm_interconnect_0:mm_to_phy_9_avalon_universal_slave_0_read -> mm_to_phy_9:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_byteenable;       // mm_interconnect_0:mm_to_phy_9_avalon_universal_slave_0_byteenable -> mm_to_phy_9:uav_byteenable
	wire         mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_readdatavalid;    // mm_to_phy_9:uav_readdatavalid -> mm_interconnect_0:mm_to_phy_9_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_lock;             // mm_interconnect_0:mm_to_phy_9_avalon_universal_slave_0_lock -> mm_to_phy_9:uav_lock
	wire         mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_write;            // mm_interconnect_0:mm_to_phy_9_avalon_universal_slave_0_write -> mm_to_phy_9:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_writedata;        // mm_interconnect_0:mm_to_phy_9_avalon_universal_slave_0_writedata -> mm_to_phy_9:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_burstcount;       // mm_interconnect_0:mm_to_phy_9_avalon_universal_slave_0_burstcount -> mm_to_phy_9:uav_burstcount
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_readdata;        // rx_sc_fifo_9:uav_readdata -> mm_interconnect_0:rx_sc_fifo_9_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_waitrequest;     // rx_sc_fifo_9:uav_waitrequest -> mm_interconnect_0:rx_sc_fifo_9_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:rx_sc_fifo_9_avalon_universal_slave_0_debugaccess -> rx_sc_fifo_9:uav_debugaccess
	wire   [4:0] mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_address;         // mm_interconnect_0:rx_sc_fifo_9_avalon_universal_slave_0_address -> rx_sc_fifo_9:uav_address
	wire         mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_read;            // mm_interconnect_0:rx_sc_fifo_9_avalon_universal_slave_0_read -> rx_sc_fifo_9:uav_read
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:rx_sc_fifo_9_avalon_universal_slave_0_byteenable -> rx_sc_fifo_9:uav_byteenable
	wire         mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_readdatavalid;   // rx_sc_fifo_9:uav_readdatavalid -> mm_interconnect_0:rx_sc_fifo_9_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_lock;            // mm_interconnect_0:rx_sc_fifo_9_avalon_universal_slave_0_lock -> rx_sc_fifo_9:uav_lock
	wire         mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_write;           // mm_interconnect_0:rx_sc_fifo_9_avalon_universal_slave_0_write -> rx_sc_fifo_9:uav_write
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_writedata;       // mm_interconnect_0:rx_sc_fifo_9_avalon_universal_slave_0_writedata -> rx_sc_fifo_9:uav_writedata
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:rx_sc_fifo_9_avalon_universal_slave_0_burstcount -> rx_sc_fifo_9:uav_burstcount
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_readdata;        // tx_sc_fifo_9:uav_readdata -> mm_interconnect_0:tx_sc_fifo_9_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_waitrequest;     // tx_sc_fifo_9:uav_waitrequest -> mm_interconnect_0:tx_sc_fifo_9_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:tx_sc_fifo_9_avalon_universal_slave_0_debugaccess -> tx_sc_fifo_9:uav_debugaccess
	wire   [4:0] mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_address;         // mm_interconnect_0:tx_sc_fifo_9_avalon_universal_slave_0_address -> tx_sc_fifo_9:uav_address
	wire         mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_read;            // mm_interconnect_0:tx_sc_fifo_9_avalon_universal_slave_0_read -> tx_sc_fifo_9:uav_read
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:tx_sc_fifo_9_avalon_universal_slave_0_byteenable -> tx_sc_fifo_9:uav_byteenable
	wire         mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_readdatavalid;   // tx_sc_fifo_9:uav_readdatavalid -> mm_interconnect_0:tx_sc_fifo_9_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_lock;            // mm_interconnect_0:tx_sc_fifo_9_avalon_universal_slave_0_lock -> tx_sc_fifo_9:uav_lock
	wire         mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_write;           // mm_interconnect_0:tx_sc_fifo_9_avalon_universal_slave_0_write -> tx_sc_fifo_9:uav_write
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_writedata;       // mm_interconnect_0:tx_sc_fifo_9_avalon_universal_slave_0_writedata -> tx_sc_fifo_9:uav_writedata
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:tx_sc_fifo_9_avalon_universal_slave_0_burstcount -> tx_sc_fifo_9:uav_burstcount
	wire  [31:0] mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_readdata;       // eth_gen_mon_9:uav_readdata -> mm_interconnect_0:eth_gen_mon_9_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_waitrequest;    // eth_gen_mon_9:uav_waitrequest -> mm_interconnect_0:eth_gen_mon_9_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:eth_gen_mon_9_avalon_universal_slave_0_debugaccess -> eth_gen_mon_9:uav_debugaccess
	wire  [13:0] mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_address;        // mm_interconnect_0:eth_gen_mon_9_avalon_universal_slave_0_address -> eth_gen_mon_9:uav_address
	wire         mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_read;           // mm_interconnect_0:eth_gen_mon_9_avalon_universal_slave_0_read -> eth_gen_mon_9:uav_read
	wire   [3:0] mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:eth_gen_mon_9_avalon_universal_slave_0_byteenable -> eth_gen_mon_9:uav_byteenable
	wire         mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_readdatavalid;  // eth_gen_mon_9:uav_readdatavalid -> mm_interconnect_0:eth_gen_mon_9_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_lock;           // mm_interconnect_0:eth_gen_mon_9_avalon_universal_slave_0_lock -> eth_gen_mon_9:uav_lock
	wire         mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_write;          // mm_interconnect_0:eth_gen_mon_9_avalon_universal_slave_0_write -> eth_gen_mon_9:uav_write
	wire  [31:0] mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_writedata;      // mm_interconnect_0:eth_gen_mon_9_avalon_universal_slave_0_writedata -> eth_gen_mon_9:uav_writedata
	wire   [3:0] mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:eth_gen_mon_9_avalon_universal_slave_0_burstcount -> eth_gen_mon_9:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_readdata;        // mm_to_mac_10:uav_readdata -> mm_interconnect_0:mm_to_mac_10_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_waitrequest;     // mm_to_mac_10:uav_waitrequest -> mm_interconnect_0:mm_to_mac_10_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:mm_to_mac_10_avalon_universal_slave_0_debugaccess -> mm_to_mac_10:uav_debugaccess
	wire  [14:0] mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_address;         // mm_interconnect_0:mm_to_mac_10_avalon_universal_slave_0_address -> mm_to_mac_10:uav_address
	wire         mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_read;            // mm_interconnect_0:mm_to_mac_10_avalon_universal_slave_0_read -> mm_to_mac_10:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:mm_to_mac_10_avalon_universal_slave_0_byteenable -> mm_to_mac_10:uav_byteenable
	wire         mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_readdatavalid;   // mm_to_mac_10:uav_readdatavalid -> mm_interconnect_0:mm_to_mac_10_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_lock;            // mm_interconnect_0:mm_to_mac_10_avalon_universal_slave_0_lock -> mm_to_mac_10:uav_lock
	wire         mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_write;           // mm_interconnect_0:mm_to_mac_10_avalon_universal_slave_0_write -> mm_to_mac_10:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_writedata;       // mm_interconnect_0:mm_to_mac_10_avalon_universal_slave_0_writedata -> mm_to_mac_10:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:mm_to_mac_10_avalon_universal_slave_0_burstcount -> mm_to_mac_10:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_readdata;        // mm_to_phy_10:uav_readdata -> mm_interconnect_0:mm_to_phy_10_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_waitrequest;     // mm_to_phy_10:uav_waitrequest -> mm_interconnect_0:mm_to_phy_10_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:mm_to_phy_10_avalon_universal_slave_0_debugaccess -> mm_to_phy_10:uav_debugaccess
	wire  [12:0] mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_address;         // mm_interconnect_0:mm_to_phy_10_avalon_universal_slave_0_address -> mm_to_phy_10:uav_address
	wire         mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_read;            // mm_interconnect_0:mm_to_phy_10_avalon_universal_slave_0_read -> mm_to_phy_10:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:mm_to_phy_10_avalon_universal_slave_0_byteenable -> mm_to_phy_10:uav_byteenable
	wire         mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_readdatavalid;   // mm_to_phy_10:uav_readdatavalid -> mm_interconnect_0:mm_to_phy_10_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_lock;            // mm_interconnect_0:mm_to_phy_10_avalon_universal_slave_0_lock -> mm_to_phy_10:uav_lock
	wire         mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_write;           // mm_interconnect_0:mm_to_phy_10_avalon_universal_slave_0_write -> mm_to_phy_10:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_writedata;       // mm_interconnect_0:mm_to_phy_10_avalon_universal_slave_0_writedata -> mm_to_phy_10:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:mm_to_phy_10_avalon_universal_slave_0_burstcount -> mm_to_phy_10:uav_burstcount
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_readdata;       // rx_sc_fifo_10:uav_readdata -> mm_interconnect_0:rx_sc_fifo_10_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_waitrequest;    // rx_sc_fifo_10:uav_waitrequest -> mm_interconnect_0:rx_sc_fifo_10_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:rx_sc_fifo_10_avalon_universal_slave_0_debugaccess -> rx_sc_fifo_10:uav_debugaccess
	wire   [4:0] mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_address;        // mm_interconnect_0:rx_sc_fifo_10_avalon_universal_slave_0_address -> rx_sc_fifo_10:uav_address
	wire         mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_read;           // mm_interconnect_0:rx_sc_fifo_10_avalon_universal_slave_0_read -> rx_sc_fifo_10:uav_read
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:rx_sc_fifo_10_avalon_universal_slave_0_byteenable -> rx_sc_fifo_10:uav_byteenable
	wire         mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_readdatavalid;  // rx_sc_fifo_10:uav_readdatavalid -> mm_interconnect_0:rx_sc_fifo_10_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_lock;           // mm_interconnect_0:rx_sc_fifo_10_avalon_universal_slave_0_lock -> rx_sc_fifo_10:uav_lock
	wire         mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_write;          // mm_interconnect_0:rx_sc_fifo_10_avalon_universal_slave_0_write -> rx_sc_fifo_10:uav_write
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_writedata;      // mm_interconnect_0:rx_sc_fifo_10_avalon_universal_slave_0_writedata -> rx_sc_fifo_10:uav_writedata
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:rx_sc_fifo_10_avalon_universal_slave_0_burstcount -> rx_sc_fifo_10:uav_burstcount
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_readdata;       // tx_sc_fifo_10:uav_readdata -> mm_interconnect_0:tx_sc_fifo_10_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_waitrequest;    // tx_sc_fifo_10:uav_waitrequest -> mm_interconnect_0:tx_sc_fifo_10_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:tx_sc_fifo_10_avalon_universal_slave_0_debugaccess -> tx_sc_fifo_10:uav_debugaccess
	wire   [4:0] mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_address;        // mm_interconnect_0:tx_sc_fifo_10_avalon_universal_slave_0_address -> tx_sc_fifo_10:uav_address
	wire         mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_read;           // mm_interconnect_0:tx_sc_fifo_10_avalon_universal_slave_0_read -> tx_sc_fifo_10:uav_read
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:tx_sc_fifo_10_avalon_universal_slave_0_byteenable -> tx_sc_fifo_10:uav_byteenable
	wire         mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_readdatavalid;  // tx_sc_fifo_10:uav_readdatavalid -> mm_interconnect_0:tx_sc_fifo_10_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_lock;           // mm_interconnect_0:tx_sc_fifo_10_avalon_universal_slave_0_lock -> tx_sc_fifo_10:uav_lock
	wire         mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_write;          // mm_interconnect_0:tx_sc_fifo_10_avalon_universal_slave_0_write -> tx_sc_fifo_10:uav_write
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_writedata;      // mm_interconnect_0:tx_sc_fifo_10_avalon_universal_slave_0_writedata -> tx_sc_fifo_10:uav_writedata
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:tx_sc_fifo_10_avalon_universal_slave_0_burstcount -> tx_sc_fifo_10:uav_burstcount
	wire  [31:0] mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_readdata;      // eth_gen_mon_10:uav_readdata -> mm_interconnect_0:eth_gen_mon_10_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_waitrequest;   // eth_gen_mon_10:uav_waitrequest -> mm_interconnect_0:eth_gen_mon_10_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_debugaccess;   // mm_interconnect_0:eth_gen_mon_10_avalon_universal_slave_0_debugaccess -> eth_gen_mon_10:uav_debugaccess
	wire  [13:0] mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_address;       // mm_interconnect_0:eth_gen_mon_10_avalon_universal_slave_0_address -> eth_gen_mon_10:uav_address
	wire         mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_read;          // mm_interconnect_0:eth_gen_mon_10_avalon_universal_slave_0_read -> eth_gen_mon_10:uav_read
	wire   [3:0] mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_byteenable;    // mm_interconnect_0:eth_gen_mon_10_avalon_universal_slave_0_byteenable -> eth_gen_mon_10:uav_byteenable
	wire         mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_readdatavalid; // eth_gen_mon_10:uav_readdatavalid -> mm_interconnect_0:eth_gen_mon_10_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_lock;          // mm_interconnect_0:eth_gen_mon_10_avalon_universal_slave_0_lock -> eth_gen_mon_10:uav_lock
	wire         mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_write;         // mm_interconnect_0:eth_gen_mon_10_avalon_universal_slave_0_write -> eth_gen_mon_10:uav_write
	wire  [31:0] mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_writedata;     // mm_interconnect_0:eth_gen_mon_10_avalon_universal_slave_0_writedata -> eth_gen_mon_10:uav_writedata
	wire   [3:0] mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_burstcount;    // mm_interconnect_0:eth_gen_mon_10_avalon_universal_slave_0_burstcount -> eth_gen_mon_10:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_readdata;        // mm_to_mac_11:uav_readdata -> mm_interconnect_0:mm_to_mac_11_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_waitrequest;     // mm_to_mac_11:uav_waitrequest -> mm_interconnect_0:mm_to_mac_11_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:mm_to_mac_11_avalon_universal_slave_0_debugaccess -> mm_to_mac_11:uav_debugaccess
	wire  [14:0] mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_address;         // mm_interconnect_0:mm_to_mac_11_avalon_universal_slave_0_address -> mm_to_mac_11:uav_address
	wire         mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_read;            // mm_interconnect_0:mm_to_mac_11_avalon_universal_slave_0_read -> mm_to_mac_11:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:mm_to_mac_11_avalon_universal_slave_0_byteenable -> mm_to_mac_11:uav_byteenable
	wire         mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_readdatavalid;   // mm_to_mac_11:uav_readdatavalid -> mm_interconnect_0:mm_to_mac_11_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_lock;            // mm_interconnect_0:mm_to_mac_11_avalon_universal_slave_0_lock -> mm_to_mac_11:uav_lock
	wire         mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_write;           // mm_interconnect_0:mm_to_mac_11_avalon_universal_slave_0_write -> mm_to_mac_11:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_writedata;       // mm_interconnect_0:mm_to_mac_11_avalon_universal_slave_0_writedata -> mm_to_mac_11:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:mm_to_mac_11_avalon_universal_slave_0_burstcount -> mm_to_mac_11:uav_burstcount
	wire  [31:0] mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_readdata;        // mm_to_phy_11:uav_readdata -> mm_interconnect_0:mm_to_phy_11_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_waitrequest;     // mm_to_phy_11:uav_waitrequest -> mm_interconnect_0:mm_to_phy_11_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_debugaccess;     // mm_interconnect_0:mm_to_phy_11_avalon_universal_slave_0_debugaccess -> mm_to_phy_11:uav_debugaccess
	wire  [12:0] mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_address;         // mm_interconnect_0:mm_to_phy_11_avalon_universal_slave_0_address -> mm_to_phy_11:uav_address
	wire         mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_read;            // mm_interconnect_0:mm_to_phy_11_avalon_universal_slave_0_read -> mm_to_phy_11:uav_read
	wire   [3:0] mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_byteenable;      // mm_interconnect_0:mm_to_phy_11_avalon_universal_slave_0_byteenable -> mm_to_phy_11:uav_byteenable
	wire         mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_readdatavalid;   // mm_to_phy_11:uav_readdatavalid -> mm_interconnect_0:mm_to_phy_11_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_lock;            // mm_interconnect_0:mm_to_phy_11_avalon_universal_slave_0_lock -> mm_to_phy_11:uav_lock
	wire         mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_write;           // mm_interconnect_0:mm_to_phy_11_avalon_universal_slave_0_write -> mm_to_phy_11:uav_write
	wire  [31:0] mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_writedata;       // mm_interconnect_0:mm_to_phy_11_avalon_universal_slave_0_writedata -> mm_to_phy_11:uav_writedata
	wire   [3:0] mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_burstcount;      // mm_interconnect_0:mm_to_phy_11_avalon_universal_slave_0_burstcount -> mm_to_phy_11:uav_burstcount
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_readdata;       // rx_sc_fifo_11:uav_readdata -> mm_interconnect_0:rx_sc_fifo_11_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_waitrequest;    // rx_sc_fifo_11:uav_waitrequest -> mm_interconnect_0:rx_sc_fifo_11_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:rx_sc_fifo_11_avalon_universal_slave_0_debugaccess -> rx_sc_fifo_11:uav_debugaccess
	wire   [4:0] mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_address;        // mm_interconnect_0:rx_sc_fifo_11_avalon_universal_slave_0_address -> rx_sc_fifo_11:uav_address
	wire         mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_read;           // mm_interconnect_0:rx_sc_fifo_11_avalon_universal_slave_0_read -> rx_sc_fifo_11:uav_read
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:rx_sc_fifo_11_avalon_universal_slave_0_byteenable -> rx_sc_fifo_11:uav_byteenable
	wire         mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_readdatavalid;  // rx_sc_fifo_11:uav_readdatavalid -> mm_interconnect_0:rx_sc_fifo_11_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_lock;           // mm_interconnect_0:rx_sc_fifo_11_avalon_universal_slave_0_lock -> rx_sc_fifo_11:uav_lock
	wire         mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_write;          // mm_interconnect_0:rx_sc_fifo_11_avalon_universal_slave_0_write -> rx_sc_fifo_11:uav_write
	wire  [31:0] mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_writedata;      // mm_interconnect_0:rx_sc_fifo_11_avalon_universal_slave_0_writedata -> rx_sc_fifo_11:uav_writedata
	wire   [3:0] mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:rx_sc_fifo_11_avalon_universal_slave_0_burstcount -> rx_sc_fifo_11:uav_burstcount
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_readdata;       // tx_sc_fifo_11:uav_readdata -> mm_interconnect_0:tx_sc_fifo_11_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_waitrequest;    // tx_sc_fifo_11:uav_waitrequest -> mm_interconnect_0:tx_sc_fifo_11_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_debugaccess;    // mm_interconnect_0:tx_sc_fifo_11_avalon_universal_slave_0_debugaccess -> tx_sc_fifo_11:uav_debugaccess
	wire   [4:0] mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_address;        // mm_interconnect_0:tx_sc_fifo_11_avalon_universal_slave_0_address -> tx_sc_fifo_11:uav_address
	wire         mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_read;           // mm_interconnect_0:tx_sc_fifo_11_avalon_universal_slave_0_read -> tx_sc_fifo_11:uav_read
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_byteenable;     // mm_interconnect_0:tx_sc_fifo_11_avalon_universal_slave_0_byteenable -> tx_sc_fifo_11:uav_byteenable
	wire         mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_readdatavalid;  // tx_sc_fifo_11:uav_readdatavalid -> mm_interconnect_0:tx_sc_fifo_11_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_lock;           // mm_interconnect_0:tx_sc_fifo_11_avalon_universal_slave_0_lock -> tx_sc_fifo_11:uav_lock
	wire         mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_write;          // mm_interconnect_0:tx_sc_fifo_11_avalon_universal_slave_0_write -> tx_sc_fifo_11:uav_write
	wire  [31:0] mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_writedata;      // mm_interconnect_0:tx_sc_fifo_11_avalon_universal_slave_0_writedata -> tx_sc_fifo_11:uav_writedata
	wire   [3:0] mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_burstcount;     // mm_interconnect_0:tx_sc_fifo_11_avalon_universal_slave_0_burstcount -> tx_sc_fifo_11:uav_burstcount
	wire  [31:0] mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_readdata;      // eth_gen_mon_11:uav_readdata -> mm_interconnect_0:eth_gen_mon_11_avalon_universal_slave_0_readdata
	wire         mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_waitrequest;   // eth_gen_mon_11:uav_waitrequest -> mm_interconnect_0:eth_gen_mon_11_avalon_universal_slave_0_waitrequest
	wire         mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_debugaccess;   // mm_interconnect_0:eth_gen_mon_11_avalon_universal_slave_0_debugaccess -> eth_gen_mon_11:uav_debugaccess
	wire  [13:0] mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_address;       // mm_interconnect_0:eth_gen_mon_11_avalon_universal_slave_0_address -> eth_gen_mon_11:uav_address
	wire         mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_read;          // mm_interconnect_0:eth_gen_mon_11_avalon_universal_slave_0_read -> eth_gen_mon_11:uav_read
	wire   [3:0] mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_byteenable;    // mm_interconnect_0:eth_gen_mon_11_avalon_universal_slave_0_byteenable -> eth_gen_mon_11:uav_byteenable
	wire         mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_readdatavalid; // eth_gen_mon_11:uav_readdatavalid -> mm_interconnect_0:eth_gen_mon_11_avalon_universal_slave_0_readdatavalid
	wire         mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_lock;          // mm_interconnect_0:eth_gen_mon_11_avalon_universal_slave_0_lock -> eth_gen_mon_11:uav_lock
	wire         mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_write;         // mm_interconnect_0:eth_gen_mon_11_avalon_universal_slave_0_write -> eth_gen_mon_11:uav_write
	wire  [31:0] mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_writedata;     // mm_interconnect_0:eth_gen_mon_11_avalon_universal_slave_0_writedata -> eth_gen_mon_11:uav_writedata
	wire   [3:0] mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_burstcount;    // mm_interconnect_0:eth_gen_mon_11_avalon_universal_slave_0_burstcount -> eth_gen_mon_11:uav_burstcount
	wire         rst_controller_reset_out_reset;                                          // rst_controller:reset_out -> [eth_gen_mon_0:reset, eth_gen_mon_10:reset, eth_gen_mon_11:reset, eth_gen_mon_1:reset, eth_gen_mon_2:reset, eth_gen_mon_3:reset, eth_gen_mon_4:reset, eth_gen_mon_5:reset, eth_gen_mon_6:reset, eth_gen_mon_7:reset, eth_gen_mon_8:reset, eth_gen_mon_9:reset, mm_interconnect_0:tx_sc_fifo_0_reset_reset_bridge_in_reset_reset, rx_sc_fifo_0:reset, rx_sc_fifo_10:reset, rx_sc_fifo_11:reset, rx_sc_fifo_1:reset, rx_sc_fifo_2:reset, rx_sc_fifo_3:reset, rx_sc_fifo_4:reset, rx_sc_fifo_5:reset, rx_sc_fifo_6:reset, rx_sc_fifo_7:reset, rx_sc_fifo_8:reset, rx_sc_fifo_9:reset, tx_sc_fifo_0:reset, tx_sc_fifo_10:reset, tx_sc_fifo_11:reset, tx_sc_fifo_1:reset, tx_sc_fifo_2:reset, tx_sc_fifo_3:reset, tx_sc_fifo_4:reset, tx_sc_fifo_5:reset, tx_sc_fifo_6:reset, tx_sc_fifo_7:reset, tx_sc_fifo_8:reset, tx_sc_fifo_9:reset]
	wire         tx_xcvr_half_clk_clk_reset_reset;                                        // tx_xcvr_half_clk:reset_n_out -> rst_controller:reset_in0

	address_decode_clk_csr clk_csr (
		.clk_out     (clk_csr_clk_clk),         //  output,  width = 1,          clk.clk
		.in_clk      (clk_csr_clk),             //   input,  width = 1,       clk_in.clk
		.reset_n     (csr_reset_n),             //   input,  width = 1, clk_in_reset.reset_n
		.reset_n_out (clk_csr_clk_reset_reset)  //  output,  width = 1,    clk_reset.reset_n
	);

	address_decode_eth_gen_mon eth_gen_mon_0 (
		.av_address        (eth_gen_mon_0_avalon_anti_slave_0_address),                              //  output,  width = 12,      avalon_anti_slave_0.address
		.av_write          (eth_gen_mon_0_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (eth_gen_mon_0_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (eth_gen_mon_0_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (eth_gen_mon_0_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.av_waitrequest    (eth_gen_mon_0_avalon_anti_slave_0_waitrequest),                          //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_eth_gen_mon eth_gen_mon_1 (
		.av_address        (eth_gen_mon_1_avalon_anti_slave_0_address),                              //  output,  width = 12,      avalon_anti_slave_0.address
		.av_write          (eth_gen_mon_1_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (eth_gen_mon_1_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (eth_gen_mon_1_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (eth_gen_mon_1_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.av_waitrequest    (eth_gen_mon_1_avalon_anti_slave_0_waitrequest),                          //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_eth_gen_mon eth_gen_mon_10 (
		.av_address        (eth_gen_mon_10_avalon_anti_slave_0_address),                              //  output,  width = 12,      avalon_anti_slave_0.address
		.av_write          (eth_gen_mon_10_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (eth_gen_mon_10_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (eth_gen_mon_10_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (eth_gen_mon_10_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.av_waitrequest    (eth_gen_mon_10_avalon_anti_slave_0_waitrequest),                          //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                                //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                           //   input,   width = 1,                    reset.reset
	);

	address_decode_eth_gen_mon eth_gen_mon_11 (
		.av_address        (eth_gen_mon_11_avalon_anti_slave_0_address),                              //  output,  width = 12,      avalon_anti_slave_0.address
		.av_write          (eth_gen_mon_11_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (eth_gen_mon_11_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (eth_gen_mon_11_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (eth_gen_mon_11_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.av_waitrequest    (eth_gen_mon_11_avalon_anti_slave_0_waitrequest),                          //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                                //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                           //   input,   width = 1,                    reset.reset
	);

	address_decode_eth_gen_mon eth_gen_mon_2 (
		.av_address        (eth_gen_mon_2_avalon_anti_slave_0_address),                              //  output,  width = 12,      avalon_anti_slave_0.address
		.av_write          (eth_gen_mon_2_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (eth_gen_mon_2_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (eth_gen_mon_2_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (eth_gen_mon_2_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.av_waitrequest    (eth_gen_mon_2_avalon_anti_slave_0_waitrequest),                          //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_eth_gen_mon eth_gen_mon_3 (
		.av_address        (eth_gen_mon_3_avalon_anti_slave_0_address),                              //  output,  width = 12,      avalon_anti_slave_0.address
		.av_write          (eth_gen_mon_3_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (eth_gen_mon_3_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (eth_gen_mon_3_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (eth_gen_mon_3_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.av_waitrequest    (eth_gen_mon_3_avalon_anti_slave_0_waitrequest),                          //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_eth_gen_mon eth_gen_mon_4 (
		.av_address        (eth_gen_mon_4_avalon_anti_slave_0_address),                              //  output,  width = 12,      avalon_anti_slave_0.address
		.av_write          (eth_gen_mon_4_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (eth_gen_mon_4_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (eth_gen_mon_4_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (eth_gen_mon_4_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.av_waitrequest    (eth_gen_mon_4_avalon_anti_slave_0_waitrequest),                          //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_eth_gen_mon eth_gen_mon_5 (
		.av_address        (eth_gen_mon_5_avalon_anti_slave_0_address),                              //  output,  width = 12,      avalon_anti_slave_0.address
		.av_write          (eth_gen_mon_5_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (eth_gen_mon_5_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (eth_gen_mon_5_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (eth_gen_mon_5_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.av_waitrequest    (eth_gen_mon_5_avalon_anti_slave_0_waitrequest),                          //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_eth_gen_mon eth_gen_mon_6 (
		.av_address        (eth_gen_mon_6_avalon_anti_slave_0_address),                              //  output,  width = 12,      avalon_anti_slave_0.address
		.av_write          (eth_gen_mon_6_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (eth_gen_mon_6_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (eth_gen_mon_6_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (eth_gen_mon_6_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.av_waitrequest    (eth_gen_mon_6_avalon_anti_slave_0_waitrequest),                          //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_eth_gen_mon eth_gen_mon_7 (
		.av_address        (eth_gen_mon_7_avalon_anti_slave_0_address),                              //  output,  width = 12,      avalon_anti_slave_0.address
		.av_write          (eth_gen_mon_7_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (eth_gen_mon_7_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (eth_gen_mon_7_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (eth_gen_mon_7_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.av_waitrequest    (eth_gen_mon_7_avalon_anti_slave_0_waitrequest),                          //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_eth_gen_mon eth_gen_mon_8 (
		.av_address        (eth_gen_mon_8_avalon_anti_slave_0_address),                              //  output,  width = 12,      avalon_anti_slave_0.address
		.av_write          (eth_gen_mon_8_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (eth_gen_mon_8_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (eth_gen_mon_8_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (eth_gen_mon_8_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.av_waitrequest    (eth_gen_mon_8_avalon_anti_slave_0_waitrequest),                          //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_eth_gen_mon eth_gen_mon_9 (
		.av_address        (eth_gen_mon_9_avalon_anti_slave_0_address),                              //  output,  width = 12,      avalon_anti_slave_0.address
		.av_write          (eth_gen_mon_9_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (eth_gen_mon_9_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (eth_gen_mon_9_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (eth_gen_mon_9_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.av_waitrequest    (eth_gen_mon_9_avalon_anti_slave_0_waitrequest),                          //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_address),       //   input,  width = 14, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_master_0 master_0 (
		.clk_clk              (clk_csr_clk_clk),               //   input,   width = 1,          clk.clk
		.clk_reset_reset      (~clk_csr_clk_reset_reset),      //   input,   width = 1,    clk_reset.reset
		.master_address       (master_0_master_address),       //  output,  width = 32,       master.address
		.master_readdata      (master_0_master_readdata),      //   input,  width = 32,             .readdata
		.master_read          (master_0_master_read),          //  output,   width = 1,             .read
		.master_write         (master_0_master_write),         //  output,   width = 1,             .write
		.master_writedata     (master_0_master_writedata),     //  output,  width = 32,             .writedata
		.master_waitrequest   (master_0_master_waitrequest),   //   input,   width = 1,             .waitrequest
		.master_readdatavalid (master_0_master_readdatavalid), //   input,   width = 1,             .readdatavalid
		.master_byteenable    (master_0_master_byteenable),    //  output,   width = 4,             .byteenable
		.master_reset_reset   ()                               //  output,   width = 1, master_reset.reset
	);

	address_decode_merlin_master_translator_0 merlin_master_translator_0 (
		.av_address        (merlin_master_translator_0_avalon_anti_master_0_address),            //   input,  width = 16,      avalon_anti_master_0.address
		.av_waitrequest    (merlin_master_translator_0_avalon_anti_master_0_waitrequest),        //  output,   width = 1,                          .waitrequest
		.av_read           (merlin_master_translator_0_avalon_anti_master_0_read),               //   input,   width = 1,                          .read
		.av_readdata       (merlin_master_translator_0_avalon_anti_master_0_readdata),           //  output,  width = 32,                          .readdata
		.av_write          (merlin_master_translator_0_avalon_anti_master_0_write),              //   input,   width = 1,                          .write
		.av_writedata      (merlin_master_translator_0_avalon_anti_master_0_writedata),          //   input,  width = 32,                          .writedata
		.uav_address       (merlin_master_translator_0_avalon_universal_master_0_address),       //  output,  width = 32, avalon_universal_master_0.address
		.uav_burstcount    (merlin_master_translator_0_avalon_universal_master_0_burstcount),    //  output,  width = 10,                          .burstcount
		.uav_read          (merlin_master_translator_0_avalon_universal_master_0_read),          //  output,   width = 1,                          .read
		.uav_write         (merlin_master_translator_0_avalon_universal_master_0_write),         //  output,   width = 1,                          .write
		.uav_waitrequest   (merlin_master_translator_0_avalon_universal_master_0_waitrequest),   //   input,   width = 1,                          .waitrequest
		.uav_readdatavalid (merlin_master_translator_0_avalon_universal_master_0_readdatavalid), //   input,   width = 1,                          .readdatavalid
		.uav_byteenable    (merlin_master_translator_0_avalon_universal_master_0_byteenable),    //  output,   width = 4,                          .byteenable
		.uav_readdata      (merlin_master_translator_0_avalon_universal_master_0_readdata),      //   input,  width = 32,                          .readdata
		.uav_writedata     (merlin_master_translator_0_avalon_universal_master_0_writedata),     //  output,  width = 32,                          .writedata
		.uav_lock          (merlin_master_translator_0_avalon_universal_master_0_lock),          //  output,   width = 1,                          .lock
		.uav_debugaccess   (merlin_master_translator_0_avalon_universal_master_0_debugaccess),   //  output,   width = 1,                          .debugaccess
		.clk               (clk_csr_clk_clk),                                                    //   input,   width = 1,                       clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                            //   input,   width = 1,                     reset.reset
	);

	address_decode_mm_to_mac mm_to_mac_0 (
		.av_address        (mac_0_avalon_anti_slave_0_address),                                    //  output,  width = 13,      avalon_anti_slave_0.address
		.av_write          (mac_0_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (mac_0_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (mac_0_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (mac_0_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (mac_0_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_address),       //   input,  width = 15, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_mac mm_to_mac_1 (
		.av_address        (mac_1_avalon_anti_slave_0_address),                                    //  output,  width = 13,      avalon_anti_slave_0.address
		.av_write          (mac_1_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (mac_1_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (mac_1_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (mac_1_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (mac_1_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_address),       //   input,  width = 15, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_mac mm_to_mac_10 (
		.av_address        (mac_10_avalon_anti_slave_0_address),                                    //  output,  width = 13,      avalon_anti_slave_0.address
		.av_write          (mac_10_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (mac_10_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (mac_10_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (mac_10_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (mac_10_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_address),       //   input,  width = 15, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                       //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                               //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_mac mm_to_mac_11 (
		.av_address        (mac_11_avalon_anti_slave_0_address),                                    //  output,  width = 13,      avalon_anti_slave_0.address
		.av_write          (mac_11_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (mac_11_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (mac_11_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (mac_11_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (mac_11_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_address),       //   input,  width = 15, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                       //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                               //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_mac mm_to_mac_2 (
		.av_address        (mac_2_avalon_anti_slave_0_address),                                    //  output,  width = 13,      avalon_anti_slave_0.address
		.av_write          (mac_2_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (mac_2_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (mac_2_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (mac_2_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (mac_2_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_address),       //   input,  width = 15, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_mac mm_to_mac_3 (
		.av_address        (mac_3_avalon_anti_slave_0_address),                                    //  output,  width = 13,      avalon_anti_slave_0.address
		.av_write          (mac_3_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (mac_3_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (mac_3_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (mac_3_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (mac_3_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_address),       //   input,  width = 15, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_mac mm_to_mac_4 (
		.av_address        (mac_4_avalon_anti_slave_0_address),                                    //  output,  width = 13,      avalon_anti_slave_0.address
		.av_write          (mac_4_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (mac_4_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (mac_4_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (mac_4_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (mac_4_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_address),       //   input,  width = 15, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_mac mm_to_mac_5 (
		.av_address        (mac_5_avalon_anti_slave_0_address),                                    //  output,  width = 13,      avalon_anti_slave_0.address
		.av_write          (mac_5_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (mac_5_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (mac_5_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (mac_5_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (mac_5_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_address),       //   input,  width = 15, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_mac mm_to_mac_6 (
		.av_address        (mac_6_avalon_anti_slave_0_address),                                    //  output,  width = 13,      avalon_anti_slave_0.address
		.av_write          (mac_6_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (mac_6_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (mac_6_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (mac_6_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (mac_6_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_address),       //   input,  width = 15, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_mac mm_to_mac_7 (
		.av_address        (mac_7_avalon_anti_slave_0_address),                                    //  output,  width = 13,      avalon_anti_slave_0.address
		.av_write          (mac_7_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (mac_7_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (mac_7_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (mac_7_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (mac_7_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_address),       //   input,  width = 15, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_mac mm_to_mac_8 (
		.av_address        (mac_8_avalon_anti_slave_0_address),                                    //  output,  width = 13,      avalon_anti_slave_0.address
		.av_write          (mac_8_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (mac_8_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (mac_8_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (mac_8_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (mac_8_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_address),       //   input,  width = 15, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_mac mm_to_mac_9 (
		.av_address        (mac_9_avalon_anti_slave_0_address),                                    //  output,  width = 13,      avalon_anti_slave_0.address
		.av_write          (mac_9_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (mac_9_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (mac_9_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (mac_9_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (mac_9_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_address),       //   input,  width = 15, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_phy mm_to_phy_0 (
		.av_address        (phy_0_avalon_anti_slave_0_address),                                    //  output,  width = 11,      avalon_anti_slave_0.address
		.av_write          (phy_0_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (phy_0_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (phy_0_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (phy_0_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (phy_0_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_address),       //   input,  width = 13, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_phy mm_to_phy_1 (
		.av_address        (phy_1_avalon_anti_slave_0_address),                                    //  output,  width = 11,      avalon_anti_slave_0.address
		.av_write          (phy_1_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (phy_1_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (phy_1_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (phy_1_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (phy_1_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_address),       //   input,  width = 13, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_phy mm_to_phy_10 (
		.av_address        (phy_10_avalon_anti_slave_0_address),                                    //  output,  width = 11,      avalon_anti_slave_0.address
		.av_write          (phy_10_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (phy_10_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (phy_10_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (phy_10_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (phy_10_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_address),       //   input,  width = 13, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                       //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                               //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_phy mm_to_phy_11 (
		.av_address        (phy_11_avalon_anti_slave_0_address),                                    //  output,  width = 11,      avalon_anti_slave_0.address
		.av_write          (phy_11_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (phy_11_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (phy_11_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (phy_11_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (phy_11_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_address),       //   input,  width = 13, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                       //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                               //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_phy mm_to_phy_2 (
		.av_address        (phy_2_avalon_anti_slave_0_address),                                    //  output,  width = 11,      avalon_anti_slave_0.address
		.av_write          (phy_2_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (phy_2_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (phy_2_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (phy_2_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (phy_2_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_address),       //   input,  width = 13, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_phy mm_to_phy_3 (
		.av_address        (phy_3_avalon_anti_slave_0_address),                                    //  output,  width = 11,      avalon_anti_slave_0.address
		.av_write          (phy_3_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (phy_3_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (phy_3_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (phy_3_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (phy_3_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_address),       //   input,  width = 13, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_phy mm_to_phy_4 (
		.av_address        (phy_4_avalon_anti_slave_0_address),                                    //  output,  width = 11,      avalon_anti_slave_0.address
		.av_write          (phy_4_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (phy_4_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (phy_4_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (phy_4_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (phy_4_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_address),       //   input,  width = 13, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_phy mm_to_phy_5 (
		.av_address        (phy_5_avalon_anti_slave_0_address),                                    //  output,  width = 11,      avalon_anti_slave_0.address
		.av_write          (phy_5_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (phy_5_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (phy_5_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (phy_5_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (phy_5_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_address),       //   input,  width = 13, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_phy mm_to_phy_6 (
		.av_address        (phy_6_avalon_anti_slave_0_address),                                    //  output,  width = 11,      avalon_anti_slave_0.address
		.av_write          (phy_6_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (phy_6_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (phy_6_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (phy_6_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (phy_6_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_address),       //   input,  width = 13, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_phy mm_to_phy_7 (
		.av_address        (phy_7_avalon_anti_slave_0_address),                                    //  output,  width = 11,      avalon_anti_slave_0.address
		.av_write          (phy_7_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (phy_7_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (phy_7_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (phy_7_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (phy_7_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_address),       //   input,  width = 13, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_phy mm_to_phy_8 (
		.av_address        (phy_8_avalon_anti_slave_0_address),                                    //  output,  width = 11,      avalon_anti_slave_0.address
		.av_write          (phy_8_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (phy_8_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (phy_8_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (phy_8_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (phy_8_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_address),       //   input,  width = 13, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_mm_to_phy mm_to_phy_9 (
		.av_address        (phy_9_avalon_anti_slave_0_address),                                    //  output,  width = 11,      avalon_anti_slave_0.address
		.av_write          (phy_9_avalon_anti_slave_0_write),                                      //  output,   width = 1,                         .write
		.av_read           (phy_9_avalon_anti_slave_0_read),                                       //  output,   width = 1,                         .read
		.av_readdata       (phy_9_avalon_anti_slave_0_readdata),                                   //   input,  width = 32,                         .readdata
		.av_writedata      (phy_9_avalon_anti_slave_0_writedata),                                  //  output,  width = 32,                         .writedata
		.av_waitrequest    (phy_9_avalon_anti_slave_0_waitrequest),                                //   input,   width = 1,                         .waitrequest
		.uav_address       (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_address),       //   input,  width = 13, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (clk_csr_clk_clk),                                                      //   input,   width = 1,                      clk.clk
		.reset             (~clk_csr_clk_reset_reset)                                              //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_sc_fifo rx_sc_fifo_0 (
		.av_address        (rx_sc_fifo_0_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (rx_sc_fifo_0_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (rx_sc_fifo_0_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (rx_sc_fifo_0_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (rx_sc_fifo_0_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_sc_fifo rx_sc_fifo_1 (
		.av_address        (rx_sc_fifo_1_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (rx_sc_fifo_1_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (rx_sc_fifo_1_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (rx_sc_fifo_1_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (rx_sc_fifo_1_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_sc_fifo rx_sc_fifo_10 (
		.av_address        (rx_sc_fifo_10_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (rx_sc_fifo_10_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (rx_sc_fifo_10_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (rx_sc_fifo_10_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (rx_sc_fifo_10_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_sc_fifo rx_sc_fifo_11 (
		.av_address        (rx_sc_fifo_11_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (rx_sc_fifo_11_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (rx_sc_fifo_11_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (rx_sc_fifo_11_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (rx_sc_fifo_11_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_sc_fifo rx_sc_fifo_2 (
		.av_address        (rx_sc_fifo_2_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (rx_sc_fifo_2_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (rx_sc_fifo_2_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (rx_sc_fifo_2_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (rx_sc_fifo_2_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_sc_fifo rx_sc_fifo_3 (
		.av_address        (rx_sc_fifo_3_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (rx_sc_fifo_3_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (rx_sc_fifo_3_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (rx_sc_fifo_3_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (rx_sc_fifo_3_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_sc_fifo rx_sc_fifo_4 (
		.av_address        (rx_sc_fifo_4_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (rx_sc_fifo_4_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (rx_sc_fifo_4_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (rx_sc_fifo_4_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (rx_sc_fifo_4_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_sc_fifo rx_sc_fifo_5 (
		.av_address        (rx_sc_fifo_5_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (rx_sc_fifo_5_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (rx_sc_fifo_5_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (rx_sc_fifo_5_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (rx_sc_fifo_5_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_sc_fifo rx_sc_fifo_6 (
		.av_address        (rx_sc_fifo_6_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (rx_sc_fifo_6_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (rx_sc_fifo_6_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (rx_sc_fifo_6_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (rx_sc_fifo_6_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_sc_fifo rx_sc_fifo_7 (
		.av_address        (rx_sc_fifo_7_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (rx_sc_fifo_7_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (rx_sc_fifo_7_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (rx_sc_fifo_7_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (rx_sc_fifo_7_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_sc_fifo rx_sc_fifo_8 (
		.av_address        (rx_sc_fifo_8_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (rx_sc_fifo_8_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (rx_sc_fifo_8_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (rx_sc_fifo_8_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (rx_sc_fifo_8_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_sc_fifo rx_sc_fifo_9 (
		.av_address        (rx_sc_fifo_9_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (rx_sc_fifo_9_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (rx_sc_fifo_9_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (rx_sc_fifo_9_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (rx_sc_fifo_9_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_rx_xcvr_clk rx_xcvr_clk (
		.clk_out     (),                    //  output,  width = 1,          clk.clk
		.in_clk      (rx_xcvr_clk_clk),     //   input,  width = 1,       clk_in.clk
		.reset_n     (sync_rx_rst_reset_n), //   input,  width = 1, clk_in_reset.reset_n
		.reset_n_out ()                     //  output,  width = 1,    clk_reset.reset_n
	);

	address_decode_tx_sc_fifo tx_sc_fifo_0 (
		.av_address        (tx_sc_fifo_0_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (tx_sc_fifo_0_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (tx_sc_fifo_0_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (tx_sc_fifo_0_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (tx_sc_fifo_0_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_tx_sc_fifo tx_sc_fifo_1 (
		.av_address        (tx_sc_fifo_1_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (tx_sc_fifo_1_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (tx_sc_fifo_1_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (tx_sc_fifo_1_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (tx_sc_fifo_1_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_tx_sc_fifo tx_sc_fifo_10 (
		.av_address        (tx_sc_fifo_10_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (tx_sc_fifo_10_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (tx_sc_fifo_10_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (tx_sc_fifo_10_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (tx_sc_fifo_10_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_tx_sc_fifo tx_sc_fifo_11 (
		.av_address        (tx_sc_fifo_11_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (tx_sc_fifo_11_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (tx_sc_fifo_11_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (tx_sc_fifo_11_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (tx_sc_fifo_11_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                               //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                          //   input,   width = 1,                    reset.reset
	);

	address_decode_tx_sc_fifo tx_sc_fifo_2 (
		.av_address        (tx_sc_fifo_2_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (tx_sc_fifo_2_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (tx_sc_fifo_2_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (tx_sc_fifo_2_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (tx_sc_fifo_2_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_tx_sc_fifo tx_sc_fifo_3 (
		.av_address        (tx_sc_fifo_3_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (tx_sc_fifo_3_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (tx_sc_fifo_3_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (tx_sc_fifo_3_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (tx_sc_fifo_3_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_tx_sc_fifo tx_sc_fifo_4 (
		.av_address        (tx_sc_fifo_4_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (tx_sc_fifo_4_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (tx_sc_fifo_4_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (tx_sc_fifo_4_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (tx_sc_fifo_4_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_tx_sc_fifo tx_sc_fifo_5 (
		.av_address        (tx_sc_fifo_5_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (tx_sc_fifo_5_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (tx_sc_fifo_5_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (tx_sc_fifo_5_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (tx_sc_fifo_5_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_tx_sc_fifo tx_sc_fifo_6 (
		.av_address        (tx_sc_fifo_6_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (tx_sc_fifo_6_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (tx_sc_fifo_6_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (tx_sc_fifo_6_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (tx_sc_fifo_6_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_tx_sc_fifo tx_sc_fifo_7 (
		.av_address        (tx_sc_fifo_7_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (tx_sc_fifo_7_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (tx_sc_fifo_7_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (tx_sc_fifo_7_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (tx_sc_fifo_7_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_tx_sc_fifo tx_sc_fifo_8 (
		.av_address        (tx_sc_fifo_8_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (tx_sc_fifo_8_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (tx_sc_fifo_8_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (tx_sc_fifo_8_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (tx_sc_fifo_8_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_tx_sc_fifo tx_sc_fifo_9 (
		.av_address        (tx_sc_fifo_9_avalon_anti_slave_0_address),                              //  output,   width = 3,      avalon_anti_slave_0.address
		.av_write          (tx_sc_fifo_9_avalon_anti_slave_0_write),                                //  output,   width = 1,                         .write
		.av_read           (tx_sc_fifo_9_avalon_anti_slave_0_read),                                 //  output,   width = 1,                         .read
		.av_readdata       (tx_sc_fifo_9_avalon_anti_slave_0_readdata),                             //   input,  width = 32,                         .readdata
		.av_writedata      (tx_sc_fifo_9_avalon_anti_slave_0_writedata),                            //  output,  width = 32,                         .writedata
		.uav_address       (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_address),       //   input,   width = 5, avalon_universal_slave_0.address
		.uav_burstcount    (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_burstcount),    //   input,   width = 4,                         .burstcount
		.uav_read          (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_read),          //   input,   width = 1,                         .read
		.uav_write         (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_write),         //   input,   width = 1,                         .write
		.uav_waitrequest   (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_waitrequest),   //  output,   width = 1,                         .waitrequest
		.uav_readdatavalid (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_readdatavalid), //  output,   width = 1,                         .readdatavalid
		.uav_byteenable    (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_byteenable),    //   input,   width = 4,                         .byteenable
		.uav_readdata      (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_readdata),      //  output,  width = 32,                         .readdata
		.uav_writedata     (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_writedata),     //   input,  width = 32,                         .writedata
		.uav_lock          (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_lock),          //   input,   width = 1,                         .lock
		.uav_debugaccess   (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_debugaccess),   //   input,   width = 1,                         .debugaccess
		.clk               (tx_xcvr_half_clk_clk_clk),                                              //   input,   width = 1,                      clk.clk
		.reset             (rst_controller_reset_out_reset)                                         //   input,   width = 1,                    reset.reset
	);

	address_decode_tx_xcvr_clk tx_xcvr_clk (
		.clk_out     (),                    //  output,  width = 1,          clk.clk
		.in_clk      (tx_xcvr_clk_clk),     //   input,  width = 1,       clk_in.clk
		.reset_n     (sync_tx_rst_reset_n), //   input,  width = 1, clk_in_reset.reset_n
		.reset_n_out ()                     //  output,  width = 1,    clk_reset.reset_n
	);

	address_decode_tx_xcvr_half_clk tx_xcvr_half_clk (
		.clk_out     (tx_xcvr_half_clk_clk_clk),         //  output,  width = 1,          clk.clk
		.in_clk      (tx_xcvr_half_clk_clk),             //   input,  width = 1,       clk_in.clk
		.reset_n     (sync_tx_half_rst_reset_n),         //   input,  width = 1, clk_in_reset.reset_n
		.reset_n_out (tx_xcvr_half_clk_clk_reset_reset)  //  output,  width = 1,    clk_reset.reset_n
	);

	address_decode_altera_mm_interconnect_181_egdbf5q mm_interconnect_0 (
		.merlin_master_translator_0_avalon_universal_master_0_address       (merlin_master_translator_0_avalon_universal_master_0_address),            //   input,  width = 32,   merlin_master_translator_0_avalon_universal_master_0.address
		.merlin_master_translator_0_avalon_universal_master_0_waitrequest   (merlin_master_translator_0_avalon_universal_master_0_waitrequest),        //  output,   width = 1,                                                       .waitrequest
		.merlin_master_translator_0_avalon_universal_master_0_burstcount    (merlin_master_translator_0_avalon_universal_master_0_burstcount),         //   input,  width = 10,                                                       .burstcount
		.merlin_master_translator_0_avalon_universal_master_0_byteenable    (merlin_master_translator_0_avalon_universal_master_0_byteenable),         //   input,   width = 4,                                                       .byteenable
		.merlin_master_translator_0_avalon_universal_master_0_read          (merlin_master_translator_0_avalon_universal_master_0_read),               //   input,   width = 1,                                                       .read
		.merlin_master_translator_0_avalon_universal_master_0_readdata      (merlin_master_translator_0_avalon_universal_master_0_readdata),           //  output,  width = 32,                                                       .readdata
		.merlin_master_translator_0_avalon_universal_master_0_readdatavalid (merlin_master_translator_0_avalon_universal_master_0_readdatavalid),      //  output,   width = 1,                                                       .readdatavalid
		.merlin_master_translator_0_avalon_universal_master_0_write         (merlin_master_translator_0_avalon_universal_master_0_write),              //   input,   width = 1,                                                       .write
		.merlin_master_translator_0_avalon_universal_master_0_writedata     (merlin_master_translator_0_avalon_universal_master_0_writedata),          //   input,  width = 32,                                                       .writedata
		.merlin_master_translator_0_avalon_universal_master_0_lock          (merlin_master_translator_0_avalon_universal_master_0_lock),               //   input,   width = 1,                                                       .lock
		.merlin_master_translator_0_avalon_universal_master_0_debugaccess   (merlin_master_translator_0_avalon_universal_master_0_debugaccess),        //   input,   width = 1,                                                       .debugaccess
		.master_0_master_address                                            (master_0_master_address),                                                 //   input,  width = 32,                                        master_0_master.address
		.master_0_master_waitrequest                                        (master_0_master_waitrequest),                                             //  output,   width = 1,                                                       .waitrequest
		.master_0_master_byteenable                                         (master_0_master_byteenable),                                              //   input,   width = 4,                                                       .byteenable
		.master_0_master_read                                               (master_0_master_read),                                                    //   input,   width = 1,                                                       .read
		.master_0_master_readdata                                           (master_0_master_readdata),                                                //  output,  width = 32,                                                       .readdata
		.master_0_master_readdatavalid                                      (master_0_master_readdatavalid),                                           //  output,   width = 1,                                                       .readdatavalid
		.master_0_master_write                                              (master_0_master_write),                                                   //   input,   width = 1,                                                       .write
		.master_0_master_writedata                                          (master_0_master_writedata),                                               //   input,  width = 32,                                                       .writedata
		.mm_to_mac_0_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_address),          //  output,  width = 15,                   mm_to_mac_0_avalon_universal_slave_0.address
		.mm_to_mac_0_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_mac_0_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_mac_0_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_mac_0_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_mac_0_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_mac_0_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_mac_0_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_mac_0_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_mac_0_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_mac_0_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_mac_0_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.mm_to_phy_0_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_address),          //  output,  width = 13,                   mm_to_phy_0_avalon_universal_slave_0.address
		.mm_to_phy_0_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_phy_0_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_phy_0_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_phy_0_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_phy_0_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_phy_0_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_phy_0_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_phy_0_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_phy_0_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_phy_0_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_phy_0_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.tx_sc_fifo_0_avalon_universal_slave_0_address                      (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_address),         //  output,   width = 5,                  tx_sc_fifo_0_avalon_universal_slave_0.address
		.tx_sc_fifo_0_avalon_universal_slave_0_write                        (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.tx_sc_fifo_0_avalon_universal_slave_0_read                         (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.tx_sc_fifo_0_avalon_universal_slave_0_readdata                     (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.tx_sc_fifo_0_avalon_universal_slave_0_writedata                    (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.tx_sc_fifo_0_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.tx_sc_fifo_0_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.tx_sc_fifo_0_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.tx_sc_fifo_0_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.tx_sc_fifo_0_avalon_universal_slave_0_lock                         (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.tx_sc_fifo_0_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_tx_sc_fifo_0_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.rx_sc_fifo_0_avalon_universal_slave_0_address                      (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_address),         //  output,   width = 5,                  rx_sc_fifo_0_avalon_universal_slave_0.address
		.rx_sc_fifo_0_avalon_universal_slave_0_write                        (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.rx_sc_fifo_0_avalon_universal_slave_0_read                         (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.rx_sc_fifo_0_avalon_universal_slave_0_readdata                     (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.rx_sc_fifo_0_avalon_universal_slave_0_writedata                    (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.rx_sc_fifo_0_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.rx_sc_fifo_0_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.rx_sc_fifo_0_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.rx_sc_fifo_0_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.rx_sc_fifo_0_avalon_universal_slave_0_lock                         (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.rx_sc_fifo_0_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_rx_sc_fifo_0_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.eth_gen_mon_0_avalon_universal_slave_0_address                     (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_address),        //  output,  width = 14,                 eth_gen_mon_0_avalon_universal_slave_0.address
		.eth_gen_mon_0_avalon_universal_slave_0_write                       (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.eth_gen_mon_0_avalon_universal_slave_0_read                        (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.eth_gen_mon_0_avalon_universal_slave_0_readdata                    (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.eth_gen_mon_0_avalon_universal_slave_0_writedata                   (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.eth_gen_mon_0_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.eth_gen_mon_0_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.eth_gen_mon_0_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.eth_gen_mon_0_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.eth_gen_mon_0_avalon_universal_slave_0_lock                        (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.eth_gen_mon_0_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_eth_gen_mon_0_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.mm_to_mac_1_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_address),          //  output,  width = 15,                   mm_to_mac_1_avalon_universal_slave_0.address
		.mm_to_mac_1_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_mac_1_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_mac_1_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_mac_1_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_mac_1_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_mac_1_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_mac_1_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_mac_1_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_mac_1_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_mac_1_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_mac_1_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.mm_to_phy_1_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_address),          //  output,  width = 13,                   mm_to_phy_1_avalon_universal_slave_0.address
		.mm_to_phy_1_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_phy_1_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_phy_1_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_phy_1_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_phy_1_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_phy_1_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_phy_1_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_phy_1_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_phy_1_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_phy_1_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_phy_1_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.rx_sc_fifo_1_avalon_universal_slave_0_address                      (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_address),         //  output,   width = 5,                  rx_sc_fifo_1_avalon_universal_slave_0.address
		.rx_sc_fifo_1_avalon_universal_slave_0_write                        (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.rx_sc_fifo_1_avalon_universal_slave_0_read                         (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.rx_sc_fifo_1_avalon_universal_slave_0_readdata                     (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.rx_sc_fifo_1_avalon_universal_slave_0_writedata                    (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.rx_sc_fifo_1_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.rx_sc_fifo_1_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.rx_sc_fifo_1_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.rx_sc_fifo_1_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.rx_sc_fifo_1_avalon_universal_slave_0_lock                         (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.rx_sc_fifo_1_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_rx_sc_fifo_1_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.tx_sc_fifo_1_avalon_universal_slave_0_address                      (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_address),         //  output,   width = 5,                  tx_sc_fifo_1_avalon_universal_slave_0.address
		.tx_sc_fifo_1_avalon_universal_slave_0_write                        (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.tx_sc_fifo_1_avalon_universal_slave_0_read                         (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.tx_sc_fifo_1_avalon_universal_slave_0_readdata                     (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.tx_sc_fifo_1_avalon_universal_slave_0_writedata                    (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.tx_sc_fifo_1_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.tx_sc_fifo_1_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.tx_sc_fifo_1_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.tx_sc_fifo_1_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.tx_sc_fifo_1_avalon_universal_slave_0_lock                         (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.tx_sc_fifo_1_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_tx_sc_fifo_1_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.eth_gen_mon_1_avalon_universal_slave_0_address                     (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_address),        //  output,  width = 14,                 eth_gen_mon_1_avalon_universal_slave_0.address
		.eth_gen_mon_1_avalon_universal_slave_0_write                       (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.eth_gen_mon_1_avalon_universal_slave_0_read                        (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.eth_gen_mon_1_avalon_universal_slave_0_readdata                    (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.eth_gen_mon_1_avalon_universal_slave_0_writedata                   (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.eth_gen_mon_1_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.eth_gen_mon_1_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.eth_gen_mon_1_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.eth_gen_mon_1_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.eth_gen_mon_1_avalon_universal_slave_0_lock                        (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.eth_gen_mon_1_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_eth_gen_mon_1_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.mm_to_mac_2_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_address),          //  output,  width = 15,                   mm_to_mac_2_avalon_universal_slave_0.address
		.mm_to_mac_2_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_mac_2_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_mac_2_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_mac_2_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_mac_2_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_mac_2_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_mac_2_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_mac_2_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_mac_2_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_mac_2_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_mac_2_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.mm_to_phy_2_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_address),          //  output,  width = 13,                   mm_to_phy_2_avalon_universal_slave_0.address
		.mm_to_phy_2_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_phy_2_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_phy_2_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_phy_2_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_phy_2_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_phy_2_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_phy_2_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_phy_2_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_phy_2_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_phy_2_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_phy_2_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.rx_sc_fifo_2_avalon_universal_slave_0_address                      (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_address),         //  output,   width = 5,                  rx_sc_fifo_2_avalon_universal_slave_0.address
		.rx_sc_fifo_2_avalon_universal_slave_0_write                        (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.rx_sc_fifo_2_avalon_universal_slave_0_read                         (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.rx_sc_fifo_2_avalon_universal_slave_0_readdata                     (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.rx_sc_fifo_2_avalon_universal_slave_0_writedata                    (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.rx_sc_fifo_2_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.rx_sc_fifo_2_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.rx_sc_fifo_2_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.rx_sc_fifo_2_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.rx_sc_fifo_2_avalon_universal_slave_0_lock                         (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.rx_sc_fifo_2_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_rx_sc_fifo_2_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.tx_sc_fifo_2_avalon_universal_slave_0_address                      (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_address),         //  output,   width = 5,                  tx_sc_fifo_2_avalon_universal_slave_0.address
		.tx_sc_fifo_2_avalon_universal_slave_0_write                        (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.tx_sc_fifo_2_avalon_universal_slave_0_read                         (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.tx_sc_fifo_2_avalon_universal_slave_0_readdata                     (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.tx_sc_fifo_2_avalon_universal_slave_0_writedata                    (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.tx_sc_fifo_2_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.tx_sc_fifo_2_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.tx_sc_fifo_2_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.tx_sc_fifo_2_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.tx_sc_fifo_2_avalon_universal_slave_0_lock                         (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.tx_sc_fifo_2_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_tx_sc_fifo_2_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.eth_gen_mon_2_avalon_universal_slave_0_address                     (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_address),        //  output,  width = 14,                 eth_gen_mon_2_avalon_universal_slave_0.address
		.eth_gen_mon_2_avalon_universal_slave_0_write                       (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.eth_gen_mon_2_avalon_universal_slave_0_read                        (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.eth_gen_mon_2_avalon_universal_slave_0_readdata                    (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.eth_gen_mon_2_avalon_universal_slave_0_writedata                   (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.eth_gen_mon_2_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.eth_gen_mon_2_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.eth_gen_mon_2_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.eth_gen_mon_2_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.eth_gen_mon_2_avalon_universal_slave_0_lock                        (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.eth_gen_mon_2_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_eth_gen_mon_2_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.mm_to_mac_3_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_address),          //  output,  width = 15,                   mm_to_mac_3_avalon_universal_slave_0.address
		.mm_to_mac_3_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_mac_3_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_mac_3_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_mac_3_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_mac_3_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_mac_3_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_mac_3_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_mac_3_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_mac_3_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_mac_3_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_mac_3_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.mm_to_phy_3_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_address),          //  output,  width = 13,                   mm_to_phy_3_avalon_universal_slave_0.address
		.mm_to_phy_3_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_phy_3_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_phy_3_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_phy_3_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_phy_3_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_phy_3_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_phy_3_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_phy_3_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_phy_3_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_phy_3_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_phy_3_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.rx_sc_fifo_3_avalon_universal_slave_0_address                      (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_address),         //  output,   width = 5,                  rx_sc_fifo_3_avalon_universal_slave_0.address
		.rx_sc_fifo_3_avalon_universal_slave_0_write                        (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.rx_sc_fifo_3_avalon_universal_slave_0_read                         (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.rx_sc_fifo_3_avalon_universal_slave_0_readdata                     (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.rx_sc_fifo_3_avalon_universal_slave_0_writedata                    (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.rx_sc_fifo_3_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.rx_sc_fifo_3_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.rx_sc_fifo_3_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.rx_sc_fifo_3_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.rx_sc_fifo_3_avalon_universal_slave_0_lock                         (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.rx_sc_fifo_3_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_rx_sc_fifo_3_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.tx_sc_fifo_3_avalon_universal_slave_0_address                      (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_address),         //  output,   width = 5,                  tx_sc_fifo_3_avalon_universal_slave_0.address
		.tx_sc_fifo_3_avalon_universal_slave_0_write                        (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.tx_sc_fifo_3_avalon_universal_slave_0_read                         (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.tx_sc_fifo_3_avalon_universal_slave_0_readdata                     (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.tx_sc_fifo_3_avalon_universal_slave_0_writedata                    (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.tx_sc_fifo_3_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.tx_sc_fifo_3_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.tx_sc_fifo_3_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.tx_sc_fifo_3_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.tx_sc_fifo_3_avalon_universal_slave_0_lock                         (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.tx_sc_fifo_3_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_tx_sc_fifo_3_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.eth_gen_mon_3_avalon_universal_slave_0_address                     (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_address),        //  output,  width = 14,                 eth_gen_mon_3_avalon_universal_slave_0.address
		.eth_gen_mon_3_avalon_universal_slave_0_write                       (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.eth_gen_mon_3_avalon_universal_slave_0_read                        (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.eth_gen_mon_3_avalon_universal_slave_0_readdata                    (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.eth_gen_mon_3_avalon_universal_slave_0_writedata                   (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.eth_gen_mon_3_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.eth_gen_mon_3_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.eth_gen_mon_3_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.eth_gen_mon_3_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.eth_gen_mon_3_avalon_universal_slave_0_lock                        (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.eth_gen_mon_3_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_eth_gen_mon_3_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.mm_to_mac_4_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_address),          //  output,  width = 15,                   mm_to_mac_4_avalon_universal_slave_0.address
		.mm_to_mac_4_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_mac_4_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_mac_4_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_mac_4_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_mac_4_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_mac_4_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_mac_4_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_mac_4_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_mac_4_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_mac_4_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_mac_4_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.mm_to_phy_4_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_address),          //  output,  width = 13,                   mm_to_phy_4_avalon_universal_slave_0.address
		.mm_to_phy_4_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_phy_4_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_phy_4_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_phy_4_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_phy_4_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_phy_4_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_phy_4_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_phy_4_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_phy_4_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_phy_4_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_phy_4_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.rx_sc_fifo_4_avalon_universal_slave_0_address                      (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_address),         //  output,   width = 5,                  rx_sc_fifo_4_avalon_universal_slave_0.address
		.rx_sc_fifo_4_avalon_universal_slave_0_write                        (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.rx_sc_fifo_4_avalon_universal_slave_0_read                         (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.rx_sc_fifo_4_avalon_universal_slave_0_readdata                     (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.rx_sc_fifo_4_avalon_universal_slave_0_writedata                    (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.rx_sc_fifo_4_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.rx_sc_fifo_4_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.rx_sc_fifo_4_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.rx_sc_fifo_4_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.rx_sc_fifo_4_avalon_universal_slave_0_lock                         (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.rx_sc_fifo_4_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_rx_sc_fifo_4_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.tx_sc_fifo_4_avalon_universal_slave_0_address                      (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_address),         //  output,   width = 5,                  tx_sc_fifo_4_avalon_universal_slave_0.address
		.tx_sc_fifo_4_avalon_universal_slave_0_write                        (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.tx_sc_fifo_4_avalon_universal_slave_0_read                         (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.tx_sc_fifo_4_avalon_universal_slave_0_readdata                     (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.tx_sc_fifo_4_avalon_universal_slave_0_writedata                    (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.tx_sc_fifo_4_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.tx_sc_fifo_4_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.tx_sc_fifo_4_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.tx_sc_fifo_4_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.tx_sc_fifo_4_avalon_universal_slave_0_lock                         (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.tx_sc_fifo_4_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_tx_sc_fifo_4_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.eth_gen_mon_4_avalon_universal_slave_0_address                     (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_address),        //  output,  width = 14,                 eth_gen_mon_4_avalon_universal_slave_0.address
		.eth_gen_mon_4_avalon_universal_slave_0_write                       (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.eth_gen_mon_4_avalon_universal_slave_0_read                        (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.eth_gen_mon_4_avalon_universal_slave_0_readdata                    (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.eth_gen_mon_4_avalon_universal_slave_0_writedata                   (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.eth_gen_mon_4_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.eth_gen_mon_4_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.eth_gen_mon_4_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.eth_gen_mon_4_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.eth_gen_mon_4_avalon_universal_slave_0_lock                        (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.eth_gen_mon_4_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_eth_gen_mon_4_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.mm_to_mac_5_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_address),          //  output,  width = 15,                   mm_to_mac_5_avalon_universal_slave_0.address
		.mm_to_mac_5_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_mac_5_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_mac_5_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_mac_5_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_mac_5_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_mac_5_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_mac_5_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_mac_5_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_mac_5_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_mac_5_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_mac_5_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.mm_to_phy_5_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_address),          //  output,  width = 13,                   mm_to_phy_5_avalon_universal_slave_0.address
		.mm_to_phy_5_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_phy_5_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_phy_5_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_phy_5_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_phy_5_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_phy_5_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_phy_5_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_phy_5_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_phy_5_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_phy_5_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_phy_5_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.rx_sc_fifo_5_avalon_universal_slave_0_address                      (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_address),         //  output,   width = 5,                  rx_sc_fifo_5_avalon_universal_slave_0.address
		.rx_sc_fifo_5_avalon_universal_slave_0_write                        (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.rx_sc_fifo_5_avalon_universal_slave_0_read                         (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.rx_sc_fifo_5_avalon_universal_slave_0_readdata                     (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.rx_sc_fifo_5_avalon_universal_slave_0_writedata                    (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.rx_sc_fifo_5_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.rx_sc_fifo_5_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.rx_sc_fifo_5_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.rx_sc_fifo_5_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.rx_sc_fifo_5_avalon_universal_slave_0_lock                         (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.rx_sc_fifo_5_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_rx_sc_fifo_5_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.tx_sc_fifo_5_avalon_universal_slave_0_address                      (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_address),         //  output,   width = 5,                  tx_sc_fifo_5_avalon_universal_slave_0.address
		.tx_sc_fifo_5_avalon_universal_slave_0_write                        (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.tx_sc_fifo_5_avalon_universal_slave_0_read                         (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.tx_sc_fifo_5_avalon_universal_slave_0_readdata                     (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.tx_sc_fifo_5_avalon_universal_slave_0_writedata                    (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.tx_sc_fifo_5_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.tx_sc_fifo_5_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.tx_sc_fifo_5_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.tx_sc_fifo_5_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.tx_sc_fifo_5_avalon_universal_slave_0_lock                         (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.tx_sc_fifo_5_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_tx_sc_fifo_5_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.eth_gen_mon_5_avalon_universal_slave_0_address                     (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_address),        //  output,  width = 14,                 eth_gen_mon_5_avalon_universal_slave_0.address
		.eth_gen_mon_5_avalon_universal_slave_0_write                       (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.eth_gen_mon_5_avalon_universal_slave_0_read                        (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.eth_gen_mon_5_avalon_universal_slave_0_readdata                    (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.eth_gen_mon_5_avalon_universal_slave_0_writedata                   (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.eth_gen_mon_5_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.eth_gen_mon_5_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.eth_gen_mon_5_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.eth_gen_mon_5_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.eth_gen_mon_5_avalon_universal_slave_0_lock                        (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.eth_gen_mon_5_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_eth_gen_mon_5_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.mm_to_mac_6_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_address),          //  output,  width = 15,                   mm_to_mac_6_avalon_universal_slave_0.address
		.mm_to_mac_6_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_mac_6_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_mac_6_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_mac_6_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_mac_6_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_mac_6_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_mac_6_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_mac_6_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_mac_6_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_mac_6_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_mac_6_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.mm_to_phy_6_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_address),          //  output,  width = 13,                   mm_to_phy_6_avalon_universal_slave_0.address
		.mm_to_phy_6_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_phy_6_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_phy_6_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_phy_6_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_phy_6_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_phy_6_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_phy_6_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_phy_6_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_phy_6_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_phy_6_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_phy_6_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.rx_sc_fifo_6_avalon_universal_slave_0_address                      (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_address),         //  output,   width = 5,                  rx_sc_fifo_6_avalon_universal_slave_0.address
		.rx_sc_fifo_6_avalon_universal_slave_0_write                        (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.rx_sc_fifo_6_avalon_universal_slave_0_read                         (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.rx_sc_fifo_6_avalon_universal_slave_0_readdata                     (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.rx_sc_fifo_6_avalon_universal_slave_0_writedata                    (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.rx_sc_fifo_6_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.rx_sc_fifo_6_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.rx_sc_fifo_6_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.rx_sc_fifo_6_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.rx_sc_fifo_6_avalon_universal_slave_0_lock                         (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.rx_sc_fifo_6_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_rx_sc_fifo_6_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.tx_sc_fifo_6_avalon_universal_slave_0_address                      (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_address),         //  output,   width = 5,                  tx_sc_fifo_6_avalon_universal_slave_0.address
		.tx_sc_fifo_6_avalon_universal_slave_0_write                        (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.tx_sc_fifo_6_avalon_universal_slave_0_read                         (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.tx_sc_fifo_6_avalon_universal_slave_0_readdata                     (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.tx_sc_fifo_6_avalon_universal_slave_0_writedata                    (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.tx_sc_fifo_6_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.tx_sc_fifo_6_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.tx_sc_fifo_6_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.tx_sc_fifo_6_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.tx_sc_fifo_6_avalon_universal_slave_0_lock                         (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.tx_sc_fifo_6_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_tx_sc_fifo_6_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.eth_gen_mon_6_avalon_universal_slave_0_address                     (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_address),        //  output,  width = 14,                 eth_gen_mon_6_avalon_universal_slave_0.address
		.eth_gen_mon_6_avalon_universal_slave_0_write                       (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.eth_gen_mon_6_avalon_universal_slave_0_read                        (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.eth_gen_mon_6_avalon_universal_slave_0_readdata                    (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.eth_gen_mon_6_avalon_universal_slave_0_writedata                   (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.eth_gen_mon_6_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.eth_gen_mon_6_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.eth_gen_mon_6_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.eth_gen_mon_6_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.eth_gen_mon_6_avalon_universal_slave_0_lock                        (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.eth_gen_mon_6_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_eth_gen_mon_6_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.mm_to_mac_7_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_address),          //  output,  width = 15,                   mm_to_mac_7_avalon_universal_slave_0.address
		.mm_to_mac_7_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_mac_7_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_mac_7_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_mac_7_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_mac_7_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_mac_7_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_mac_7_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_mac_7_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_mac_7_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_mac_7_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_mac_7_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.mm_to_phy_7_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_address),          //  output,  width = 13,                   mm_to_phy_7_avalon_universal_slave_0.address
		.mm_to_phy_7_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_phy_7_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_phy_7_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_phy_7_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_phy_7_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_phy_7_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_phy_7_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_phy_7_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_phy_7_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_phy_7_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_phy_7_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.rx_sc_fifo_7_avalon_universal_slave_0_address                      (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_address),         //  output,   width = 5,                  rx_sc_fifo_7_avalon_universal_slave_0.address
		.rx_sc_fifo_7_avalon_universal_slave_0_write                        (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.rx_sc_fifo_7_avalon_universal_slave_0_read                         (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.rx_sc_fifo_7_avalon_universal_slave_0_readdata                     (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.rx_sc_fifo_7_avalon_universal_slave_0_writedata                    (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.rx_sc_fifo_7_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.rx_sc_fifo_7_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.rx_sc_fifo_7_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.rx_sc_fifo_7_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.rx_sc_fifo_7_avalon_universal_slave_0_lock                         (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.rx_sc_fifo_7_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_rx_sc_fifo_7_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.tx_sc_fifo_7_avalon_universal_slave_0_address                      (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_address),         //  output,   width = 5,                  tx_sc_fifo_7_avalon_universal_slave_0.address
		.tx_sc_fifo_7_avalon_universal_slave_0_write                        (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.tx_sc_fifo_7_avalon_universal_slave_0_read                         (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.tx_sc_fifo_7_avalon_universal_slave_0_readdata                     (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.tx_sc_fifo_7_avalon_universal_slave_0_writedata                    (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.tx_sc_fifo_7_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.tx_sc_fifo_7_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.tx_sc_fifo_7_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.tx_sc_fifo_7_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.tx_sc_fifo_7_avalon_universal_slave_0_lock                         (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.tx_sc_fifo_7_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_tx_sc_fifo_7_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.eth_gen_mon_7_avalon_universal_slave_0_address                     (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_address),        //  output,  width = 14,                 eth_gen_mon_7_avalon_universal_slave_0.address
		.eth_gen_mon_7_avalon_universal_slave_0_write                       (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.eth_gen_mon_7_avalon_universal_slave_0_read                        (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.eth_gen_mon_7_avalon_universal_slave_0_readdata                    (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.eth_gen_mon_7_avalon_universal_slave_0_writedata                   (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.eth_gen_mon_7_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.eth_gen_mon_7_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.eth_gen_mon_7_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.eth_gen_mon_7_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.eth_gen_mon_7_avalon_universal_slave_0_lock                        (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.eth_gen_mon_7_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_eth_gen_mon_7_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.mm_to_mac_8_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_address),          //  output,  width = 15,                   mm_to_mac_8_avalon_universal_slave_0.address
		.mm_to_mac_8_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_mac_8_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_mac_8_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_mac_8_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_mac_8_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_mac_8_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_mac_8_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_mac_8_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_mac_8_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_mac_8_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_mac_8_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.mm_to_phy_8_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_address),          //  output,  width = 13,                   mm_to_phy_8_avalon_universal_slave_0.address
		.mm_to_phy_8_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_phy_8_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_phy_8_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_phy_8_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_phy_8_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_phy_8_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_phy_8_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_phy_8_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_phy_8_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_phy_8_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_phy_8_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.rx_sc_fifo_8_avalon_universal_slave_0_address                      (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_address),         //  output,   width = 5,                  rx_sc_fifo_8_avalon_universal_slave_0.address
		.rx_sc_fifo_8_avalon_universal_slave_0_write                        (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.rx_sc_fifo_8_avalon_universal_slave_0_read                         (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.rx_sc_fifo_8_avalon_universal_slave_0_readdata                     (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.rx_sc_fifo_8_avalon_universal_slave_0_writedata                    (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.rx_sc_fifo_8_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.rx_sc_fifo_8_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.rx_sc_fifo_8_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.rx_sc_fifo_8_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.rx_sc_fifo_8_avalon_universal_slave_0_lock                         (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.rx_sc_fifo_8_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_rx_sc_fifo_8_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.tx_sc_fifo_8_avalon_universal_slave_0_address                      (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_address),         //  output,   width = 5,                  tx_sc_fifo_8_avalon_universal_slave_0.address
		.tx_sc_fifo_8_avalon_universal_slave_0_write                        (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.tx_sc_fifo_8_avalon_universal_slave_0_read                         (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.tx_sc_fifo_8_avalon_universal_slave_0_readdata                     (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.tx_sc_fifo_8_avalon_universal_slave_0_writedata                    (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.tx_sc_fifo_8_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.tx_sc_fifo_8_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.tx_sc_fifo_8_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.tx_sc_fifo_8_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.tx_sc_fifo_8_avalon_universal_slave_0_lock                         (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.tx_sc_fifo_8_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_tx_sc_fifo_8_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.eth_gen_mon_8_avalon_universal_slave_0_address                     (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_address),        //  output,  width = 14,                 eth_gen_mon_8_avalon_universal_slave_0.address
		.eth_gen_mon_8_avalon_universal_slave_0_write                       (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.eth_gen_mon_8_avalon_universal_slave_0_read                        (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.eth_gen_mon_8_avalon_universal_slave_0_readdata                    (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.eth_gen_mon_8_avalon_universal_slave_0_writedata                   (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.eth_gen_mon_8_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.eth_gen_mon_8_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.eth_gen_mon_8_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.eth_gen_mon_8_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.eth_gen_mon_8_avalon_universal_slave_0_lock                        (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.eth_gen_mon_8_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_eth_gen_mon_8_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.mm_to_mac_9_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_address),          //  output,  width = 15,                   mm_to_mac_9_avalon_universal_slave_0.address
		.mm_to_mac_9_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_mac_9_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_mac_9_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_mac_9_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_mac_9_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_mac_9_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_mac_9_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_mac_9_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_mac_9_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_mac_9_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_mac_9_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.mm_to_phy_9_avalon_universal_slave_0_address                       (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_address),          //  output,  width = 13,                   mm_to_phy_9_avalon_universal_slave_0.address
		.mm_to_phy_9_avalon_universal_slave_0_write                         (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_write),            //  output,   width = 1,                                                       .write
		.mm_to_phy_9_avalon_universal_slave_0_read                          (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_read),             //  output,   width = 1,                                                       .read
		.mm_to_phy_9_avalon_universal_slave_0_readdata                      (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_readdata),         //   input,  width = 32,                                                       .readdata
		.mm_to_phy_9_avalon_universal_slave_0_writedata                     (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_writedata),        //  output,  width = 32,                                                       .writedata
		.mm_to_phy_9_avalon_universal_slave_0_burstcount                    (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_burstcount),       //  output,   width = 4,                                                       .burstcount
		.mm_to_phy_9_avalon_universal_slave_0_byteenable                    (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_byteenable),       //  output,   width = 4,                                                       .byteenable
		.mm_to_phy_9_avalon_universal_slave_0_readdatavalid                 (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_readdatavalid),    //   input,   width = 1,                                                       .readdatavalid
		.mm_to_phy_9_avalon_universal_slave_0_waitrequest                   (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_waitrequest),      //   input,   width = 1,                                                       .waitrequest
		.mm_to_phy_9_avalon_universal_slave_0_lock                          (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_lock),             //  output,   width = 1,                                                       .lock
		.mm_to_phy_9_avalon_universal_slave_0_debugaccess                   (mm_interconnect_0_mm_to_phy_9_avalon_universal_slave_0_debugaccess),      //  output,   width = 1,                                                       .debugaccess
		.rx_sc_fifo_9_avalon_universal_slave_0_address                      (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_address),         //  output,   width = 5,                  rx_sc_fifo_9_avalon_universal_slave_0.address
		.rx_sc_fifo_9_avalon_universal_slave_0_write                        (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.rx_sc_fifo_9_avalon_universal_slave_0_read                         (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.rx_sc_fifo_9_avalon_universal_slave_0_readdata                     (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.rx_sc_fifo_9_avalon_universal_slave_0_writedata                    (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.rx_sc_fifo_9_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.rx_sc_fifo_9_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.rx_sc_fifo_9_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.rx_sc_fifo_9_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.rx_sc_fifo_9_avalon_universal_slave_0_lock                         (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.rx_sc_fifo_9_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_rx_sc_fifo_9_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.tx_sc_fifo_9_avalon_universal_slave_0_address                      (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_address),         //  output,   width = 5,                  tx_sc_fifo_9_avalon_universal_slave_0.address
		.tx_sc_fifo_9_avalon_universal_slave_0_write                        (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.tx_sc_fifo_9_avalon_universal_slave_0_read                         (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.tx_sc_fifo_9_avalon_universal_slave_0_readdata                     (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.tx_sc_fifo_9_avalon_universal_slave_0_writedata                    (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.tx_sc_fifo_9_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.tx_sc_fifo_9_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.tx_sc_fifo_9_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.tx_sc_fifo_9_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.tx_sc_fifo_9_avalon_universal_slave_0_lock                         (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.tx_sc_fifo_9_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_tx_sc_fifo_9_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.eth_gen_mon_9_avalon_universal_slave_0_address                     (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_address),        //  output,  width = 14,                 eth_gen_mon_9_avalon_universal_slave_0.address
		.eth_gen_mon_9_avalon_universal_slave_0_write                       (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.eth_gen_mon_9_avalon_universal_slave_0_read                        (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.eth_gen_mon_9_avalon_universal_slave_0_readdata                    (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.eth_gen_mon_9_avalon_universal_slave_0_writedata                   (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.eth_gen_mon_9_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.eth_gen_mon_9_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.eth_gen_mon_9_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.eth_gen_mon_9_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.eth_gen_mon_9_avalon_universal_slave_0_lock                        (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.eth_gen_mon_9_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_eth_gen_mon_9_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.mm_to_mac_10_avalon_universal_slave_0_address                      (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_address),         //  output,  width = 15,                  mm_to_mac_10_avalon_universal_slave_0.address
		.mm_to_mac_10_avalon_universal_slave_0_write                        (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.mm_to_mac_10_avalon_universal_slave_0_read                         (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.mm_to_mac_10_avalon_universal_slave_0_readdata                     (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.mm_to_mac_10_avalon_universal_slave_0_writedata                    (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.mm_to_mac_10_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.mm_to_mac_10_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.mm_to_mac_10_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.mm_to_mac_10_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.mm_to_mac_10_avalon_universal_slave_0_lock                         (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.mm_to_mac_10_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_mm_to_mac_10_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.mm_to_phy_10_avalon_universal_slave_0_address                      (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_address),         //  output,  width = 13,                  mm_to_phy_10_avalon_universal_slave_0.address
		.mm_to_phy_10_avalon_universal_slave_0_write                        (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.mm_to_phy_10_avalon_universal_slave_0_read                         (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.mm_to_phy_10_avalon_universal_slave_0_readdata                     (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.mm_to_phy_10_avalon_universal_slave_0_writedata                    (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.mm_to_phy_10_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.mm_to_phy_10_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.mm_to_phy_10_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.mm_to_phy_10_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.mm_to_phy_10_avalon_universal_slave_0_lock                         (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.mm_to_phy_10_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_mm_to_phy_10_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.rx_sc_fifo_10_avalon_universal_slave_0_address                     (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_address),        //  output,   width = 5,                 rx_sc_fifo_10_avalon_universal_slave_0.address
		.rx_sc_fifo_10_avalon_universal_slave_0_write                       (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.rx_sc_fifo_10_avalon_universal_slave_0_read                        (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.rx_sc_fifo_10_avalon_universal_slave_0_readdata                    (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.rx_sc_fifo_10_avalon_universal_slave_0_writedata                   (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.rx_sc_fifo_10_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.rx_sc_fifo_10_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.rx_sc_fifo_10_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.rx_sc_fifo_10_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.rx_sc_fifo_10_avalon_universal_slave_0_lock                        (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.rx_sc_fifo_10_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_rx_sc_fifo_10_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.tx_sc_fifo_10_avalon_universal_slave_0_address                     (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_address),        //  output,   width = 5,                 tx_sc_fifo_10_avalon_universal_slave_0.address
		.tx_sc_fifo_10_avalon_universal_slave_0_write                       (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.tx_sc_fifo_10_avalon_universal_slave_0_read                        (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.tx_sc_fifo_10_avalon_universal_slave_0_readdata                    (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.tx_sc_fifo_10_avalon_universal_slave_0_writedata                   (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.tx_sc_fifo_10_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.tx_sc_fifo_10_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.tx_sc_fifo_10_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.tx_sc_fifo_10_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.tx_sc_fifo_10_avalon_universal_slave_0_lock                        (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.tx_sc_fifo_10_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_tx_sc_fifo_10_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.eth_gen_mon_10_avalon_universal_slave_0_address                    (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_address),       //  output,  width = 14,                eth_gen_mon_10_avalon_universal_slave_0.address
		.eth_gen_mon_10_avalon_universal_slave_0_write                      (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_write),         //  output,   width = 1,                                                       .write
		.eth_gen_mon_10_avalon_universal_slave_0_read                       (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_read),          //  output,   width = 1,                                                       .read
		.eth_gen_mon_10_avalon_universal_slave_0_readdata                   (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_readdata),      //   input,  width = 32,                                                       .readdata
		.eth_gen_mon_10_avalon_universal_slave_0_writedata                  (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_writedata),     //  output,  width = 32,                                                       .writedata
		.eth_gen_mon_10_avalon_universal_slave_0_burstcount                 (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_burstcount),    //  output,   width = 4,                                                       .burstcount
		.eth_gen_mon_10_avalon_universal_slave_0_byteenable                 (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_byteenable),    //  output,   width = 4,                                                       .byteenable
		.eth_gen_mon_10_avalon_universal_slave_0_readdatavalid              (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_readdatavalid), //   input,   width = 1,                                                       .readdatavalid
		.eth_gen_mon_10_avalon_universal_slave_0_waitrequest                (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_waitrequest),   //   input,   width = 1,                                                       .waitrequest
		.eth_gen_mon_10_avalon_universal_slave_0_lock                       (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_lock),          //  output,   width = 1,                                                       .lock
		.eth_gen_mon_10_avalon_universal_slave_0_debugaccess                (mm_interconnect_0_eth_gen_mon_10_avalon_universal_slave_0_debugaccess),   //  output,   width = 1,                                                       .debugaccess
		.mm_to_mac_11_avalon_universal_slave_0_address                      (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_address),         //  output,  width = 15,                  mm_to_mac_11_avalon_universal_slave_0.address
		.mm_to_mac_11_avalon_universal_slave_0_write                        (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.mm_to_mac_11_avalon_universal_slave_0_read                         (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.mm_to_mac_11_avalon_universal_slave_0_readdata                     (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.mm_to_mac_11_avalon_universal_slave_0_writedata                    (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.mm_to_mac_11_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.mm_to_mac_11_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.mm_to_mac_11_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.mm_to_mac_11_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.mm_to_mac_11_avalon_universal_slave_0_lock                         (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.mm_to_mac_11_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_mm_to_mac_11_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.mm_to_phy_11_avalon_universal_slave_0_address                      (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_address),         //  output,  width = 13,                  mm_to_phy_11_avalon_universal_slave_0.address
		.mm_to_phy_11_avalon_universal_slave_0_write                        (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_write),           //  output,   width = 1,                                                       .write
		.mm_to_phy_11_avalon_universal_slave_0_read                         (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_read),            //  output,   width = 1,                                                       .read
		.mm_to_phy_11_avalon_universal_slave_0_readdata                     (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_readdata),        //   input,  width = 32,                                                       .readdata
		.mm_to_phy_11_avalon_universal_slave_0_writedata                    (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_writedata),       //  output,  width = 32,                                                       .writedata
		.mm_to_phy_11_avalon_universal_slave_0_burstcount                   (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_burstcount),      //  output,   width = 4,                                                       .burstcount
		.mm_to_phy_11_avalon_universal_slave_0_byteenable                   (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_byteenable),      //  output,   width = 4,                                                       .byteenable
		.mm_to_phy_11_avalon_universal_slave_0_readdatavalid                (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_readdatavalid),   //   input,   width = 1,                                                       .readdatavalid
		.mm_to_phy_11_avalon_universal_slave_0_waitrequest                  (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_waitrequest),     //   input,   width = 1,                                                       .waitrequest
		.mm_to_phy_11_avalon_universal_slave_0_lock                         (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_lock),            //  output,   width = 1,                                                       .lock
		.mm_to_phy_11_avalon_universal_slave_0_debugaccess                  (mm_interconnect_0_mm_to_phy_11_avalon_universal_slave_0_debugaccess),     //  output,   width = 1,                                                       .debugaccess
		.rx_sc_fifo_11_avalon_universal_slave_0_address                     (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_address),        //  output,   width = 5,                 rx_sc_fifo_11_avalon_universal_slave_0.address
		.rx_sc_fifo_11_avalon_universal_slave_0_write                       (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.rx_sc_fifo_11_avalon_universal_slave_0_read                        (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.rx_sc_fifo_11_avalon_universal_slave_0_readdata                    (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.rx_sc_fifo_11_avalon_universal_slave_0_writedata                   (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.rx_sc_fifo_11_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.rx_sc_fifo_11_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.rx_sc_fifo_11_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.rx_sc_fifo_11_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.rx_sc_fifo_11_avalon_universal_slave_0_lock                        (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.rx_sc_fifo_11_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_rx_sc_fifo_11_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.tx_sc_fifo_11_avalon_universal_slave_0_address                     (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_address),        //  output,   width = 5,                 tx_sc_fifo_11_avalon_universal_slave_0.address
		.tx_sc_fifo_11_avalon_universal_slave_0_write                       (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_write),          //  output,   width = 1,                                                       .write
		.tx_sc_fifo_11_avalon_universal_slave_0_read                        (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_read),           //  output,   width = 1,                                                       .read
		.tx_sc_fifo_11_avalon_universal_slave_0_readdata                    (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_readdata),       //   input,  width = 32,                                                       .readdata
		.tx_sc_fifo_11_avalon_universal_slave_0_writedata                   (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_writedata),      //  output,  width = 32,                                                       .writedata
		.tx_sc_fifo_11_avalon_universal_slave_0_burstcount                  (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_burstcount),     //  output,   width = 4,                                                       .burstcount
		.tx_sc_fifo_11_avalon_universal_slave_0_byteenable                  (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_byteenable),     //  output,   width = 4,                                                       .byteenable
		.tx_sc_fifo_11_avalon_universal_slave_0_readdatavalid               (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_readdatavalid),  //   input,   width = 1,                                                       .readdatavalid
		.tx_sc_fifo_11_avalon_universal_slave_0_waitrequest                 (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_waitrequest),    //   input,   width = 1,                                                       .waitrequest
		.tx_sc_fifo_11_avalon_universal_slave_0_lock                        (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_lock),           //  output,   width = 1,                                                       .lock
		.tx_sc_fifo_11_avalon_universal_slave_0_debugaccess                 (mm_interconnect_0_tx_sc_fifo_11_avalon_universal_slave_0_debugaccess),    //  output,   width = 1,                                                       .debugaccess
		.eth_gen_mon_11_avalon_universal_slave_0_address                    (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_address),       //  output,  width = 14,                eth_gen_mon_11_avalon_universal_slave_0.address
		.eth_gen_mon_11_avalon_universal_slave_0_write                      (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_write),         //  output,   width = 1,                                                       .write
		.eth_gen_mon_11_avalon_universal_slave_0_read                       (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_read),          //  output,   width = 1,                                                       .read
		.eth_gen_mon_11_avalon_universal_slave_0_readdata                   (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_readdata),      //   input,  width = 32,                                                       .readdata
		.eth_gen_mon_11_avalon_universal_slave_0_writedata                  (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_writedata),     //  output,  width = 32,                                                       .writedata
		.eth_gen_mon_11_avalon_universal_slave_0_burstcount                 (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_burstcount),    //  output,   width = 4,                                                       .burstcount
		.eth_gen_mon_11_avalon_universal_slave_0_byteenable                 (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_byteenable),    //  output,   width = 4,                                                       .byteenable
		.eth_gen_mon_11_avalon_universal_slave_0_readdatavalid              (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_readdatavalid), //   input,   width = 1,                                                       .readdatavalid
		.eth_gen_mon_11_avalon_universal_slave_0_waitrequest                (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_waitrequest),   //   input,   width = 1,                                                       .waitrequest
		.eth_gen_mon_11_avalon_universal_slave_0_lock                       (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_lock),          //  output,   width = 1,                                                       .lock
		.eth_gen_mon_11_avalon_universal_slave_0_debugaccess                (mm_interconnect_0_eth_gen_mon_11_avalon_universal_slave_0_debugaccess),   //  output,   width = 1,                                                       .debugaccess
		.merlin_master_translator_0_reset_reset_bridge_in_reset_reset       (~clk_csr_clk_reset_reset),                                                //   input,   width = 1, merlin_master_translator_0_reset_reset_bridge_in_reset.reset
		.tx_sc_fifo_0_reset_reset_bridge_in_reset_reset                     (rst_controller_reset_out_reset),                                          //   input,   width = 1,               tx_sc_fifo_0_reset_reset_bridge_in_reset.reset
		.clk_csr_clk_clk                                                    (clk_csr_clk_clk),                                                         //   input,   width = 1,                                            clk_csr_clk.clk
		.tx_xcvr_half_clk_clk_clk                                           (tx_xcvr_half_clk_clk_clk)                                                 //   input,   width = 1,                                   tx_xcvr_half_clk_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~tx_xcvr_half_clk_clk_reset_reset), //   input,  width = 1, reset_in0.reset
		.clk            (tx_xcvr_half_clk_clk_clk),          //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),    //  output,  width = 1, reset_out.reset
		.reset_req      (),                                  // (terminated),                       
		.reset_req_in0  (1'b0),                              // (terminated),                       
		.reset_in1      (1'b0),                              // (terminated),                       
		.reset_req_in1  (1'b0),                              // (terminated),                       
		.reset_in2      (1'b0),                              // (terminated),                       
		.reset_req_in2  (1'b0),                              // (terminated),                       
		.reset_in3      (1'b0),                              // (terminated),                       
		.reset_req_in3  (1'b0),                              // (terminated),                       
		.reset_in4      (1'b0),                              // (terminated),                       
		.reset_req_in4  (1'b0),                              // (terminated),                       
		.reset_in5      (1'b0),                              // (terminated),                       
		.reset_req_in5  (1'b0),                              // (terminated),                       
		.reset_in6      (1'b0),                              // (terminated),                       
		.reset_req_in6  (1'b0),                              // (terminated),                       
		.reset_in7      (1'b0),                              // (terminated),                       
		.reset_req_in7  (1'b0),                              // (terminated),                       
		.reset_in8      (1'b0),                              // (terminated),                       
		.reset_req_in8  (1'b0),                              // (terminated),                       
		.reset_in9      (1'b0),                              // (terminated),                       
		.reset_req_in9  (1'b0),                              // (terminated),                       
		.reset_in10     (1'b0),                              // (terminated),                       
		.reset_req_in10 (1'b0),                              // (terminated),                       
		.reset_in11     (1'b0),                              // (terminated),                       
		.reset_req_in11 (1'b0),                              // (terminated),                       
		.reset_in12     (1'b0),                              // (terminated),                       
		.reset_req_in12 (1'b0),                              // (terminated),                       
		.reset_in13     (1'b0),                              // (terminated),                       
		.reset_req_in13 (1'b0),                              // (terminated),                       
		.reset_in14     (1'b0),                              // (terminated),                       
		.reset_req_in14 (1'b0),                              // (terminated),                       
		.reset_in15     (1'b0),                              // (terminated),                       
		.reset_req_in15 (1'b0)                               // (terminated),                       
	);

endmodule
