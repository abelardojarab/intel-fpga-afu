`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tyyv1792nCz1FyQM61+6TOFMSXmEvBZzmikDZKrAsWViqyaZuVcMeKs/Qcj83W5r
ziDRS74K/nQ7F7riP8/Fgo3nX8eM3ovZGXTewIbRWKsVEYVtOI/QOLNlWB80l4ec
1Xn3h/TtNjUUNad5JQNbaIz68UkRTAjNkBUo4lHdylo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31744)
2mfbJvacLd7Lt6loKG9pq6XL4Q0xS1KWp+1GUDCJuNR5jfBXuleqO+UTfnuOX0NJ
fMLzkYH93IUZviv8614lHiFwXEbVzO8XWIYXKqWKdUPnKwE0PWzszzUTmVhSjtaq
pBo1dxMvTof9742HO6DotPcpYCqEhqRK8+XHxB6fUZeJUmBkG+6pxYTDvUmUN0BR
7LRm1bKLypC6ADl2x4q3hJBM+UfEt9kCAkSisc0z/nWaYP4upzSUF/WdVpiJluFu
W3DMsq/dUm71bmBYatM6X6eZHckOqgvv1pKV5NUInrNmXziDpSyCPNI0QdYJN2sW
UZ6MCkDySW+WoKKegrGuj0O3rnsuOvnn4aSdW4I4Jtr2PJDrJ5jKv+STZpv9+YGG
KnUowJKiVnSPexhsiabpAZBJ+eQabYmNiqaPGmAy0DyZimuI7I2RPTULdmZ2Cken
fd5fmVldHDj8wm8UAphBuJT5XhiqIthTlf8c+JMhBsyiWlKiUb0uSve9oLOA2STz
EbIcyM7XEjiO3+4Q3sGQWzESgbMZbRRPQ2J+i821R5Uth4IVosv3oV5Ql+saE4Q6
IzU4uzZhFhk7jY2Av2lAO+6xpsUWrV5h86r2TpJu9WdwlDiYg8vJisY8QyAbnkko
Zz68q0oeLcAqaliT1MIP86L3ENrgK5mYRyn3R+5b269fSkRamMXjiBcLO5mTl7Z9
MNuAHxbTTuat8pEJ3TGCzzDGFlBePE2M7dZwLzRFQrrqDGKGwSeyfSEhdmv0ZIig
gkbrZUh2kDuL+KIdrfbiLvjuPbOJ+t9CgpoHTosNDR4tJhI32kcsOAGNXsmRbQiF
iUNhg4Dzzhtzr8291jvA2koQ8vsG4OIyqrgobK9HFA5PrwG6am/w9GgKhRY5uWW2
zHtzxfmKxQhmfdxlv5r+e/XQr8ND+thTlloP8AZihTbvkYgyas6TVANiVNwwROxV
mHPq5jAqigqRkGmMNijW4k3xCJIYG+Wd4541B6umCZoxwJi1G6jqV9+7siZIIhJ4
5655gSyP7S/JPEfY1uOJAy5APR6ImSCb3W18HVcG2M6Vgqcn/MjWEwgvnThTRoCF
qaNYw0GHY7KjMFh/VTdorgU0Fqib3XnhFRBRtAD+LyMhrA6srrX6/Pd93zx3Q7jl
N/jSMZSfOclV1BkX5727gKpz0D2ALaQwGr9EOpzmZ2MoC4hq6GBygWkjVtwU9G3Y
ChlKHK+nZEk69u9bGVJIR56hSlHxcmaSVUQiItwjYEtwgyrbjm+VNRVR7FlrojET
AAunn3ImebCozrG0V1LRL7SMmfWKsywslw5ZtaAcxAbQQlUn9FNRDNO7hW/QAlqI
GYrAG1l1pzW6WxlqnUAM2NS9DnW+pE771W8+lYhr5bG0AWD8Sbu7O52GpCuNW8ED
KyETVOs3PcJcfqmgL84WRrHjanIe0Pu3WZfMUHW5E9Pb1jUWeuy7/BfF8ENX63AL
jCDxItPbKXw3pE6U85p133XJvRk9lMiCUnkd9odHTjm7mDgCXREsaWfwNCqRzToQ
wkDh/Hlc2kmF+PwFlDupmIi/rm+c3qyR8HHXghvHGKCqZIvwiLHx4Wui2UvS7hli
D1MtTfCRQ71SqbUUBDtX7u8G/oVFVFYSQknl2jvsLLrxzkbV+j90xEczWeQuF0xf
NGpZguRdnbxgtnvXnF3MX/ly9wNrom7tcRR77XoPAPPVMY9Z4tpHl6obK36koLy7
++/eYnuBzrMr+rT+Ws5p9KDMcpdc19WfMxcAOqlNfrRwb7KngOMRiqKGCtOC8JYW
K8wzKIRBU9/bGgYtUiYVBujeG6Pd0sKfkZOlz0jVDAIZuk3lst8rVjpXzugsR9mq
k6PS7vQLcvMYuTbng5xXk2on+/uVBN+oqTTnqjfaBpkZx54TUXT6pdVmG88Pzxbc
RTKAf0n1cO+3P0Dv1C1WbOFRRi2o81xE02+Ka8ePDtsRtv33lyfiBjdt1eEs7zfq
BMaZQL5MUcPoOra0UPpTWYwkrizPMt8slUnI3QBCx2iBkDrSNROQ7Y+YD4taT6jO
rTfr7/qP92VgaVgu6lATQWLfXeny9dzfmwnzSVkOsQnbiVWJDJixbVBEksGhEpnd
6PLCEqDq60PUmDcQqnvD4z5RIAM+XgeVPSHW9UthZTmsf80lwNmJNMx/Q0vaQe7d
U1CKdRaNjzgMWoszEEXpe4sKe79kL8hTdNYJhldrjWDd5AZ6BKM5U+4qveB+wdLO
VpwAoiaooMvvUgQe2Erd/pmBIdiN8TF3VAxBBW/7zgxbOnQxnZGQwQCuchEnuI/U
7Jc6p3Qb3bWJ6Pb+wropYpH7sMKBkFMI0K5Ez3I1UFL0le8Mp7O6E+5ockFxzTnU
nPjQXVztseBwqxjKkpjw7OPR3l2Lu89yrx3A6LHJwXJ+JGbXOz5aQh9wgQNTmWSm
5ONIgazls7lj9TlZDkKtM7irdcaejaWEPsZxTCt/getiATaAPUZ85eNBWMt13JmM
RAFSM0AvQP+cxKrgmeMCyY9N1B4qIzmccmVjn4p78yP/NHhDtIPr9I1BsYgGHY3k
2Q1+KqV9rKJWjCLSVD8FaMms4mC91nRMM2vhj1K2O9d5xIXZSzU4yZDZfpOX4QyZ
xHtpnhr5vUbC97m9QL1l6xVchJsIzejZ86K2/ibLFe5yUxIFgmfjZmPVy7eA4UHU
m1Fe0jkAa8G+wv6xUwRj0Fx0xV76elf8Ql9lxRW6uSdpCidxTdpD7Ek/cmXfSdGs
6BVsA7D/iLndiV0a/QNtfF8TZYnH10fk+wICg1KkuR9FBhzTAiWMEhbKa6/Jy7sB
5TiO5lE5kOzXtXrdoMGBWcTI5n923ZTxRRIhbTpV0Lj6mtlbmGie7w8s9M84p+Yl
HKJUgJOaNCnfPmeqw9h6yqiJKbwfvGOTuqB6aNzywHDdBVDwIlA2jB6+0eTmXboM
QMsexSKGT1DqWvgQYEbaiUwDME3+bbZ6ROGxK5lGvSTC0RbW7rznisULZOoGe6yy
AZqWx1wJIk2+mv3xsLdMnNyN9xEYp8+/SBqfPApJO15bGYP3X0W4rG3rhdGydx1i
S2umV6vH6+JJGthla/RbOMRMs+otGTGcn+DsrXknUG2PhS6sCcMYsVWtcT++LQ/0
BcWq4IT+XgYDXPHRPHfuPZs9ENWvVmk6jayybWLiNao7F6u+lrWoFzSyLTn2M2uN
1tGlA68rvh89jX8Pf7pi0QmhYnJl3CBHPZmgiWq6Mx9v5LOk1SwkuwHI0uw+PlWE
xyUakgfVdOfhMocobK/9huh6ZUMV9ZBQzTS9lRi5vzieosn1gFjZnLw9YLdVD6Pt
kAZLDkkFKdDsYHnQyzFXKJT67+EN8zUyjYDWnRydyZGc+w5r9F4tvPXw7drhZ80l
qriJhjaz7aaqdYzYr9PuGkY4f5lc+D1hxQWOb8SkiJPIvqIQzQkuNcnxHUsXePFa
kfJomRtShmYs4LfaxWUCyvh41fnBI89cCabX4BqKciDU1j8lsRdzBLKXmW/LmPR0
1WzhrlvWp2Vi05DTRo2RJ9g6+zNXBb28xXToXxJlm8VlD/PNX0qiza6S11ST3Brp
gXJIisbvVCAO2sMm3NB+avJFz0pKd4w+zpwMD6k5J8mhrFYnj5880VRB7lyKr1xc
P/fF+RXOjcP6myaVXfDbHywOuLVv5kyQFeKRqIKt9cTsGFcSkEo2gKLtAhQk8INL
1R8D7ifBj2pvrSS4/pwkK6/TaZcMYNKkjJvgWa2/6e4zR0b7WgXX5CSwr8qUIfUi
6z5UAbi6/PZys95fbfvQASEa5/U2RdPiyfD2MhWGraqHnoK8tow18laT51FWnBhu
CZjNXAu0SajmphD3lUs5q2/6E1QKvBvcs97JZ9PS5e385sv5D4KheMmuukrQAuyt
U4BT8qNzhDvGFVUvr4NkKM5GTas5BLl4vWV6bDdgqEfBeI5YPwbD99aw44/FJsww
02YdvcFBfesSnp1WhcPBAtJviEmdRd/8WDrZy5zUegGQ/K5BvFgkTK5lxq1R9aUV
rlZJWs+oubMKTNFauvjjjxWK+6NpYQI8VxVeurMQlGDTQ4nY60Op0eH5LYj9erau
gHEyYddJNdAMIds0jf4bre4UJWZyrOZFztJDcyLpGe3CWgXeHYepbBTqwhEUWZp/
JhF9zI2S/3BrS2PZimqKznwUH1VTAW8J6g9lJDiLt3V1UKUaDnmu22+sAeNEOWF4
gOMrmtfteQawQ4+0Hk7e73ycjdO3m9BpYek5UpZoDf2hfxAW+ZhLplGYsXjMT6Gx
VGmRQnvgea32EQoXRsXg8yxOUeb2nskVnhMzBuOFuA1XQrAtOWsc60JewHG2Y0VQ
OAXPEXvpN8nYYmBQAoX0MpmfcOCeSANjTwrggThjTbauc3ooezBiu1EZ2b+ZHBt8
EJUGbmUTqBRxKsw/6U+mB09YGBJhhVYCkjDPE3zRWxYDgTXqNC/gsj/0nlUhJBo3
gtFn5aPtc9cLbz7M6sZdx/R35+8kKjuCiFlJx1x9kjAu9QqL1vwSnaF7Zp7/v75s
L4cXiBg54okrW+/k+FcybLTb2VTvq2e9lDtvMrzlBAAtQZUL67mf+hJSZVhurdO2
4IiiXlnFy2ntAqJcXm+JR0RRGlbntgNeFDXvmoqD5FGoTbJeVsh7OavNlFyfPbgI
FotacV7SQF5IbmUm/5VWfWJowvqaIS3H1+Swz0RX1smmyIW4zylNZIHEjp1QgPCZ
2Wn5CIhyTxgftsc+dbfo2wikieoRZMi2TPZHeUoJzLc6ocVAzSPZBEROOp4/k0B6
jnv9iQ11p4LSYf7XKXYLIEmPcMF+CmSIa4zNehYtk0FlnJK2iTrph3hRTt7Yrz7t
5z9dArF4yt4LKKlC8RCCAZsy5v7wFgkYeTJM1SODcPHgIod6TFh4zS2WdXbIJtTZ
lxCQSd/DfQLQPNmYjTqniJpgWbGXjMXOx5FfXECov0vh7f0ugyGWtMRUDzRfMYJo
M8Qh8vp6hsnu7J1x628IsLWM9f+AW0P2zv7isC+J+kZjecppxzqJpIL/ZkZ9yjwc
x0jqaGZ2soSHiHV9f32OzXkRat46+0rZJ/KlTkQZpxeNZUC9Pasmffz1w/Xn+4dc
GpjvgQfvgAN4Z+7LwgidPzX+BqhHOxZw6V2II5dnRewl5BFZ+MDtXTjUQkBgFNze
KmmTqIY7ZyzmefZvJdelm+f4/HSM1yOYz5wl67T0jJfpC89pi9So6gvUkf/Dryei
cToM4qk78jrlVjFBLCrja5TM04xHDzUjfMHEVF+yCcg4GUo/1KHFjRervZMoqjES
h7KA45eTw8y+yzl3CCvDDjFO6VVfpCK5KFlKMIG5V5JemEY0a1LvOnRQTgQWXa5l
GnjEnugiFitcjuLL5UDhyIqv7RtcyS6bDe4MYzJ0x3WEOoV8TWDLNy2cQU0K3Tpm
LmAET8N3W5h+CzjWT8nkIHdNtxoYy/2bhlHC7sMOsHJUBJDpyZgZzAtSELtHhsws
IQf0/qyX9qgs6Uhp9VixSLXDX83e2v3gaoZY33pCJ0970q70rneTOmodpZ43H7ZK
NFSLKKcdGoBqnvbLQzWpHyu+yeBi28dWzBYhhgVfKo7LEDBBRiP7m/PBObOoYatX
e6OGcqjjISg9441IKhJH2wxsPhMc5W2HTDdl5ZG8LWOY8uKNpX4QdDND7ADav2Jt
V3jrcW39rMIvfKFQGpEQUIKskV0tzMQNYAnJEbA9x2D+gnsy+c1vLRsQQSbx6gDL
mdCPhXP8cCgR8IFwvIP3MpoLIPxoJqqWQcK14YF9c6nl6YIzqpDs1eTnY/HbUBXJ
n5wbMfLpvLYiyC+A3YhH2pEMxJSGEgktd9wia6dFTrYWMi5YHkOy7luk3DXkySLq
W5xukBWRPP0OGeF/elsfhtOQlUVTTQ7kjJCLHUNpBWhThks3urezVBANP4CltzfZ
Kzwb1gO3ikbxelKSdZxSA3tmTmzJPyQPSFQSQeIi+UPzfS8TtxzZVvkxOuMuYU4g
2ky+XvwQVgXhaPTqCVvI5HWZR+Aoqykvwgfbwwmxe8S2VvetJ+m1+lR9DlLOiqhm
anLzRbfjSZCwHmczFyz41OMvfQN1dSM53N14X0aRerX9dnL0PDI9MIAfBom4Wl2F
MlF254CTv39L8BicoUR4Yh7Zk/29MkxfzMLoAsUhjgSYcsqwUxIjsjY9qDRyndip
AdI6zqzrCoa65nJ8MlvEHwjdT/juNrAwOTvuFZqNYYAHnNfucvNxVM6wkyDSD7m0
JYQ0kpXWH+lOuTEPvunERqohqkJ41IVT5eMrM15SKg1APYZmrSm0AGAnYf9bUl9s
XtKKkoqofkijF22EWagh/0VV2l50XSMMS4yFNlzZZaD+Rgbx0NdhhpK98UkyHndx
iQBJUAENxv6daA83f822cmtAI1jKdsrBLNoTTl6tD0A2q3l6UuY0tqrUu0d8spD5
0ZoIywAA2bcHH2+gwJ9bjYd5Rvj9Eoyt22iVJ4la+/OXGO/1mfs+5CoQKWgasXYP
YQpL06NPc+0jNNDxpuZttKzsWR2Gk/Zu4bzIFtZrZQ3PhsCPXIbrAbiL64jkspPK
D48rN15zMsIRrJomepQl8ZTuy4AOegg4iKpLfeSW6ai3kQmP6tnw3vW2Dev1FUR6
5jWDVCUx2AG1qxP/pO1Ctv7jQp/6kaC6x+IIik08omLufHoYxOuv8fCtMzLaynNS
cFnGwssSoBhW2wt0KNGH5QdptHweCJnAe51KJH0xNIxXzN0uPA748NNyXgSG/eDY
L0Rhfytd+wGTeZ+UJKosKcdj3h8P4MAUZZ6OMCf0myJLM4a0uhAV+f8GK7w8PH73
x2xuBm2XslJHEmlqmUYHMziCTntjle4SvXBMXXH92FYHBFMl+XQ0lqnj3Js1IJoy
CCuazW+kQWIOwaV8orbQLoZAU+o96Vo+xJ80SkaKuqqGikabF8fWO69SYQLSEusb
d7J7DOdeudXEx0jjBDIpNhdGzm+9ET5YjKRB49Nu1YCIC2djGT+GP8vb0i8o1nAP
3rg1uKuKFLLIFX8KiF4FGM/Lj7qEsrRHfMN0JQuTcSQJyheypAE2GBXDs6iv06hs
0uJW+R3nkgrbTD2LYQwQbxtI+w0kdFXCZaBWlUv9NGYKHFy0hww6xa6hsdDkcSbb
Z5phgNmEyMXKmdC2DZhviGoQqV3PuswEZz26pZcRbn7QP05CGdfovOM8Ld7EA4mR
YiWrCookdOSKuaRi0pvu6bXBdACXo/Us47jDb3GpTFMDE1E1cYisYLu0SctvCWta
UxxTYUd0vuKQtgoA9XRdt1P0Au6yzPQrOO2dBvY7SARpnWTEcEyHWIxqm6tvEaRp
J8oHL6RPIUXkNXv0poXhlUZhHyKXk1B9IPh83WtdOIXJiuDwLuy1i/f756ysxIuN
cTkucOElHzBeID3qrtpgcnmfFBBQj6v1n/JJUtANu1TpO+2wdPYqxnLhzpbsVKvb
vgvrBRxTyrnrXWY036xj2xRLdLQUUR+38kJ0DpaM+RrGqA+nKTK2bBCnxMxAM7PH
nNNCKamrNIUsAjJewhxOPkQrki3VqeO6UGafVUrkZsvZ/qDU/Ok3jksSP9dDihK9
kPm3q9aKohpfokoKcKN5rDLZ1d1sxOG72XX3HjQGtnJYPVtsGQkGxnyeYRy1na5F
+vKz/uSM8Bs1q5OG3w4z4TcLLEJWnMOPeM/5uQbntIK0XYGwunJ4W65g7+5oecLN
jinySwlxkQcVztTujYwTkRs1xv8BQBR7JQX3g3IXUMz9zp76K6xxXwJU9/Co1YVD
bB96hfmmokYl8BxTk/Q8bjzIv/IXw6Msv64oIpx/tiDu6/qqmY988gBm2embnGCH
8fQ6uUjvW8Eo4M9ppHhYiwhy7cb+uG1XRyOBGTphneNaI+yKkY7mxdH4WjgwPqxt
jhgqHX3fn1ZFJUB+w3/Bu3DzYpryCLBGawiiKgBBXycmWtaVYtsEnv5Vpm6BfP0N
9v126ytuoIKI63F8FCyOqgNKfyfetkcz+kE41/aEzqcNhxj11SXSWBInyC1D+QNX
+Uwxkajq6bVrLdhW4zjxg6sycyxDd2BR883f+z4xAn7LoLSoYVo8fUS/6tlDQvoH
g8MBENgRBAxbwHU7Kp/8wx2cNuCEOpNC8RXgoCVf+3xIaj3QsALXNG7g2bw58X9C
aq6++1dQvOaGShZJMnI4Xuo6TYOzz3wEruch3Feopz7sHZ5UsgSk7gqBLmMDL+M2
hObDvWeBv8plc/JiZHTdOHOjILhIqsNl0z5Cl1DIUr8rYiW1Rh0oon4q3B5voSAw
3DG+Z+gU+VbgXjaiCIawVmWdkQezQOf/97i8wGSBfQg/KHgsLNUGNsS5KmSy5XZL
/oJGbh7VB/4UqWQVPGrncBtM86TWQbwoRDohsd4W3yRsc8aJQXSQVuOSEYgE8J6D
8OJZBG1BmiGX+ehpoh7oNHFUjBFNDwzzYlxyFPFsNm9RnYofna/0XwrUEEAcp4zM
yr7ruBwZcGe9BAwumAbWd0G6E/TxiFDhN4QpD2LWwGgh191hCZWoitlkQdgEc/CV
iQ1qYZv22CHjtVQ8i05kqoIqeX+2VF3aZtE4aqGW3vW2LFdDHvho0OzSOYqNZDUG
wltEImmgajopIGsXcNkBQF0ZdemPqJNCdw5NtKXRLca3jfHTSw6zIDOY9E5SLjjR
eWkJ0xezgn7aPqng6WMYTn385H0LOx59+w7R8GFlQB//NPZ3THp4H0OKM3zsXAPk
I3JdHqctdx0UW9nZPie533zL351a41gX8HX4pVYuWWEejXqchGS+6Rs1IqGxaQn1
EskRr0hX/w0++cS5teWmyWBrwCld+HzQED4rmDQ9AyzXbCioU0/IcMGbtgsNX1ey
efGomqEfAfbX5/ciR1z7DA+lxt9kZjvK1ZSH2JRCrqMf8xpTepHj37e8eX2CjO46
i9iWPyo3OvxgMr1EDaMBn+wcLFgZ/cFXtFwOFtgbCYq2aRJE3v++VfDJ5fq6RKCB
sGJ76EcB9oRox0fhwStEiK3GKSo1uxz7F2Bv0faa9+0sHZLVpjjuTRng3ZOfApI6
d5vK5WDG2VzjMw5R6smWjYlIeoLmp5NaX+xteU8NG4p0x71RqXZdfDDiC7T4hDgm
7VpNEgbtuN1Ms1PlNUl7o0YPzvDBUIMeiqbMew3hEJCxbJksepheh0vOHUxPtW3a
bjDElPosunZYL2mQgrZSkfhrccRgYfSxBBfr3U7C0dLUaR+cjCg17oQbHFyInHBB
X/TuXX7jAZ6U4hrxApaINURB3gLiVp6qK0Wbm4KELXutSZNmaOVBJIyug+nm1pJp
aqEJcIs7ERAnf6MP5eQwD7rt0LoEjg4dktxkD1bVsiuTloz53P/mywqlk1LJNfMS
gcXiOArEc1tcqG0Nz+DEvrbXoDJmzUw+DcQGs/giG+arYppjxwaFo6cjnOVCN9gL
CiphECrVlf1NPsThyS0KCQLXJn0Yo+isbur4Faqz+3CuvDUsMFhedt8KG6k86Cle
0gZL0qwrZoJ1sEkZThilzhAX3Yovn4t5AXfMFSorbENww8VGSZ2PgXu19R1MyRZG
MQgj/9oSiezrZFezTvheaAy3Dxe5CvZseKK88SnOq4idl3tPFeOVqI99BoTc/6jL
NfsNYKgENLA9mvAaAx6+IqD0aqUUGcfY0MLiQAvMV/tfGR5G1egeVXNDkZ2mG2qt
K5T7jg0vAH5LAXL62XbBwH0tgjH4Ovow3O6hkOF5GepLiZ8J+9J+6vFcqYa/3aAz
BucFE6BgINPQjbEOD7MslCgYEpKhjGxYiGLRi7zW685/eusDbsWGqU3fi1iYWlem
QwIbsuAPLCOh/hU5M22JjEeaAbpmIm3IgybfsjrgqJKzM9bqPH1+je6EvABPCcwN
gvpUt8ueZnbUi/ax0fTykdV/FNje4hu6RREcouapBfJmP3gd6rgYmPkO7Jkc+vlE
Wl+NgzhsM6pZVDVsKp4BiROSbtQsOFhU+7VzM3nMOSd+FOHqKNfvPCgSTxV9NJXB
fGiPPeasdb9zKrMylAr1GKqHH3/WzThN/8ozIcw9OYu5aB1Xxee9CmnThw260yFB
mnvlu0bz+th/zmhBFSU2je9B1GUuCIpvWo26ROk6z8NNutsyu2WV3AuaiyPzGUtJ
PS9h6sZ8sSwKUcuvlwzi5vUQwVtPf6usFB+6k7MhLBvSx7/axB9ZP4k2aHXhEPJz
cRQyQYt6ZCAdqgUcAxxufKb7yIaf93c8MNDCwvaIXJh/MJkTEJxtc7/rlPUAMiV2
p3CoXiORUl1fesiGOEo0qERl6Z1+XJyDmv5+n2dCTOeecBfFEnjmh/aYMPe8tW9j
H7tUU9NFzg68CvM6sOE7SrX/TNRKq/F9XDaVf900CeKyQ41fW5WJZhM9pUwct9Iy
eghIM1yecfVJheqG3HCW9sw/whFjI+0IhgZRoTnGNmTo0+HFxyil12MCwdxGzTDP
K/VL4h8evf7+IzI3zqSr8DsHBg6WRVurTmycFdpoNZpM+VuTLb/++CNT7X2Fqi7t
IVEmVzVS0wWQYsVG9O9/uizAvjNvunn516HyG1dJdWpgz7aSK1U3Vaep0pSPtNx6
CJRJTQLe5bQOC+6EB8uuZjr3mAZf61UzGmPb6RSXspLffnAjhfKHMzln+TBklUde
sjeQ1b7ew5Sfy1VzNOgqHAX5S3hwRwgFI3G5dZVSVjE06RcTZvJp9kTueSKSnBbF
jZBtuz4r1pgCqgzg/2HnXaSxcjGI5E+NmAG2gFIuZQVeANYzJICwc0pF9nOSJoZg
nqciWLauHeywpQ6FpA+Zgu3eZHXRN1vdCcwf39NFtds+bBvN+BTSM5Gagjqn4sxT
UqDBzTSMqh+Z97zXuGU+L5JmZSCFpvkGW4QkNnuQpNl4MGffV/lQN8N8yGR17hzN
TmZe5D0MTSZYWrYdwPKIqfNhhRaa+ctSjt3riAT1jE/z0zYLs88ad0YsLfsnv1LZ
DoPyt0HmbIEJpQms87BwshlALEkirKdRmIEmP8BPy091OcPOoNI33smlP/KI5rNe
Gn0esnzPeja3aANGFZ5hoE6S5l2dl0putDV5C2nY77VRBWt+AkXp5ixv2IulY1Cl
8OuaOjHRKyDn29At54cJoqpux6WqCvKOzdakZHmLCik74JoTXc3UhwyS4fGXHZgb
vuKpXFCLEGoO+xs5YzmrWq2me2PMbztvNt1tLOl13pDB9nv895khg5Wm6c2k1vcW
K93CKUGVSWfUpEQLzlHQwM9SDZ2Hrx31dZkgsd45CLKuaZmfw230QxhGLewE8rfu
KTePRexJCIY3g3PkOKMnZ1GnZUImiTZnRJIo6juwn7h+444oF6uawGTilPCZLj8M
/wT+yoDFiKC75ckminEAr0DJ7O2yCfJdYy7fug6fC96VzQul8PaC0vCHRjXDzzzS
qdSVIIUsUeaBw8/dJfeZgwx0csUZPhntu+Ym8rIXJS1I2Z588gRkZgybwNH0VJTC
UiR4kjNPf2WwB75UzVtO7YSHRF4c6CX/8xr5DAUO8iLNTW5OBkm+/cX+iQ/SgdCX
YsmYxPAB8Rwx6LNHwvFfFA4FAtUTlN1pBjVRhK/bf1SVup+MAWPcxgTCy2LxpLd/
C1cnvdgEpValnLyQfPGvWuDwCz0KJMFEOzCYjVlVLwOgdW21P4Eglf0Ez6CAH4dU
qzKWwehA/ci4JKzh/MZ6GOXkqs8CQJXzhPiOLP4KkssAw2u/53xaKmqBildb18vD
baycaYAFcZhMSRAWsLfWyRr20uPdKOVvO2JhXtC34Fo/i5/ZRs/b73SbxLgilYh0
5+MGuUSA8HwdMxN9rJ4HSQ1T2FAHg1ydUBd5PKO7lgaF22P2CIvhPm6uK+kIQ5j9
gnyEkkawudhqF9ir5RNBEklX/tt8nTn9Y/bv6yIDX1ZBvi564S8DJsvCKCvLoI2y
cU6zLJPqG6i9ARI6RhYFnfoo75EMcQNeqeEt2t9vaZ/z787EZbCJSDHoKfJZ+iIc
HxnHye/nW1Q/RqS9MDxEJWlu3qp7vPDC8IQe/Au07Efms9sUycSEmWoMnj76Ayzy
gafQgZl2lJZapPNEkT+QkCiuJZK0BwarKSe9tQHDV/C7CPrvoBFSpz3ihv/vylUN
ugOvJ50WqCpfZwk7hADXySdufs3d2Tnx7MAP9RLXK+J4DOR4ZIUhaBtVM7wyxDSl
3bBTdCQQtFRN/2JdOCjc0dw3Eiq0RWhxZaEvpCvDxYRpU9nonSSnO1UMcGOCO8f4
d3mUkG/AccmSAdXSEnHE14tMeW6Z9ZHNe1zNmEix76SPGo1tqqMXCDeCOcIKXbGk
QEKZJ+wESMdXJYGyPgakyt5KJaa0OYk1UEw7exlqbb6wZU2VeoSZBdC9RmI81WFz
v4qtKpCbkhn+VVhGG8CNkJ8QdTjgkg5AVZw23uHDFR1JARMVW3JR+WvIDiqH8OQ8
FsJ6HHnIEzVwMuqhx1ZkDD9l1ZA+YP93bV7i2X7BvMC/8WFBVOb4zQAaCTakGsu0
9ukKcc08KBzJEkL1/3IQs8KHkSFfC6D1+S8827E0M3FlZUACqgpN9Y9s3FCOMglw
VGYal9rya6JoP+zgFLzbcno4/HCtNUpIRAYdi2ND6AEKMdurcv0NQP2Lx2e3YkxP
9qfU2VbtsQ3QtIVKKM/H9cJdrNFxXGAbyM77/0uh3EY48t0fPVMFcvCguUZv8kqa
A4HrkRYxgCZJUeOkeZG6fDUI18pRHLeLOkMAUa2rJuUhtD2agtMzADsWn9o0qpLx
OUEW7YqdbBifGJoWIGsKSuFMAe0ccAaqr9hTFUDE43DfGD6PpS8HPJWP+Y6tcYsM
zw2ronmg5IYjZm0iSQaYtnya2iA3WSNnAYxJeXo5cNnKV8OKyYI2K1W2zS9P42X7
8M5mcv3GVl4HBvZB/5A9uw/jfunw/FoJLiHvXp7Om8rdXVCQ+3vBT42ch6RYjtRq
HolW9krAv5nkwD8BHrQ5p7NNSpOzSa9WmFIFS1BJK+r+IFdiiaawKDy/TOoiqixD
wmwHPknrVdBzrt5owwbTRwL6GOgShykxs7pM4B8WzMMk7TTMgXltFT1XUnqsDS87
nsf5/RwprSmu4vF3hyOCbfTOgOR2h9WhjY5nWdGlgMX1wa/PFzq7uvJ7llZT1ulv
OeXjyvLoDJhVXoyhu7sMwAPBDoMIfDoB5J8nm5PHjrhcVZf5iihSGo5EK8apa1v3
hFJbjSEuVftOrzl5875v6k5giJLOzCwoOCDwQfQ5oDZ4LEsi/fzjHinAvu0JN/iW
VIK0w06N15YmGqFwCsXL+Ws1Z+zUdbYzdDS98TSZNB7zF99Icf2QyXWOiaaQ5YS3
VlRMzXQL13JeIhIkdGmKKhGG8xGhv952iOvWqN+/dKk8jkEj6dXs3+PMERkoN/fG
OQwIm6P7Jom6DdaXa/DQDfErqpnx5VoVi2s9wNHzD4iR/TrVSPcGVHf4RoW43MEU
GQLbIWHonyX7iVwUSF2LAcgPWAsnBZifmgTBCsf2T/Evt0EABBybK2Yzrn4CGZem
ISZ8UZhpBC5TfTzKmY0/3uwW1R0NdwzNyrAf+D9i3P6v6w47sKHgeRi8xkDCd7T0
+Q6bKH/wA48zVhzEx+N0KcFL7m6VvvE//aX2a0aS03WACIwezhXsAANMvN7DunjU
RVP+ZobF2l8YLWlJyh/E0RRytpX1XCem7K6ntGtJLL2I9QFN/wVb/ImHqEOmUFze
KOQXDkx+RoP3PbcwAgrBI/Cl2E92pV+xWm8juNjXw7rD0JcrI0VmlT2cRNEATlGR
k5QS7vBU4w91a8X+WBPakwhzpPbWXCiPZ4vqPvbbHd1FnVkxqruItFBBmw33FXA5
niLrUZR9WgHfdv1Opj6inzt8tWXj1pFHN+M8QdgChDDFJOfx2PhzlBihSmkuZ+Sp
ELaQ0wKOfpoEVQ73cakpUktWp9wP2HzN8Nx8v/8mpCAFctMriakfA605Xpdyn1KZ
vnrklTVeRVBAUBEc84Ku/dJ2/bcomAk9rmX/4+Kz4m8fzyychwhpJ4hNWWz3QNru
LqZLZ5OYIJXqMMRqcZTOd75N4IHV6OHlVJGRHjKjaxnB3O3ZLSxHdbM4VVSX2L8+
nHBoBht6PaqdkW6dZz5XkbXgj8l9Utb7NUWcD+0hphSvPWTE3cqnMAld1ZsSHzIe
/nKap6UBsw6Nv8DSfZPoIK2Y4flFkn1uMeYNlt0lA/SR0xxghT8x8T8qOi/KREjJ
Vdj+ulTPuS37lXbIX8ZvVxBzw7H7Tgcf2E1RoAn7czkopX8AfGCsroluR2rP0IXS
7RZeuq0HbSGkdKZdJPVDjWcgyHHtq9ompHpUxo7aCCT/cOtyxleUqeliXSUAkieo
BeCljqSndynfwbZdJm1Z+W2dHbEsMoa2AY3zb6XL5RJ7WxkZhWg5RUg39fVYpk4r
LXC/55HrYVLIMNULrbQKwZXf8waO9PjlvLdLZ3iixwNaBTjVpkYkB7uFwzc5NrYI
nHxAaRjFp2suQnm9BTMWYm7SRVyvmh8it216zOELvksnyHb4Mhrv0Mg+SLZ+ngSn
O37E85OfVqEkYQgRbHIaNNz9temHc/xE7arKQMkuwlqZqVgkT+MIhmayQfs9UI8L
AVoJRJiP5sRuga3e/WG4avAHySNrcxR+Fa3hCIccck6U3Q8N60IBsPEhjuZqrRJl
tZA8dZsuC5sZYsxPkA+hpungnia+XAnP7njH5sPCBVpADljrCaaKa6wYNUQlL+QI
ZGQLcogYgDy9Adxw3qaOkqIM7lhhjvU2QUI5FubtaS2bHMJRXwtrsKckOWzzFbKT
hvWmTI9tkSEnTcL2HkLBp4tEUwddQY5zTuMYbN3f8HAY1cBhWqZ5gjVDIWaK01I0
m/yZpaM5Qwtw7bko5euJ7Sv+3HMBHV/Mz2flfYb9WbIB3B5RVAXAVoQqALFXQD5e
gIolluxfTMEx/K9o2fr8bYGPhaIzgb0y558GWsoiGA7sC7Yydu8S7T0C4ggZDkaV
44zgKZY2WEGFwEA/KXxsqSQJP9QCRMsKN44nlgidsDSqJ9deFiE9vRJfwc1u4KAm
aG45e/zlTLLzc1nKpfTKVTW6dw8fccBGVqTioHq1o+Yjf8dlS3M5Pcwq6N5st51+
83VTyELbTEK3uS72ca3oyMGfaioHkHPRfGFYCkXNWUuNfQKRBxHqBKJSy0VgYT37
Qc1jDGnPgzze9mYqWkNADqiELpqVyeS8SDRoKknxkuA6bo4hcktr0lHweEDYQaqg
MzifMAygs8eHmCAFrCXSg+Wx/MFZNef12kCN5Doul9oNpv+FA7cLFSN9vsR9ZbfD
nHHhcGEEHzyZfFcWBv4Bq6Yaht5cQEnswfiV59d+eO0eBdg5RxCCNxGOH7jOi6om
u0ftaVpPWpibG3EY3jifMe2ZaOfFzZFu6V6BV5oeRWtZhN3FjKG4W/hXMOvqhvxe
NbOJRL/Pjn/sSgipsyn3LDj6b5dNYuWELQuDdjhSUh+HH/PSmQ/eOGqdCZyCPEN8
FwSyztRGBjcdlFamnXHSjR6fUcAID3IGN7aD7549CzC3Xe+Cq0LmfyysO/ydgbED
jfpYJ/apG6WdYP6mZDjRFY3PDQE+Jzdxn4GhMcVBPiH6vFDzFSyEWmIn9p1eLO6n
NqiIEkYJqvR+piGUOkuWQ/gz071D9aon+CimOLgALPcmkKkEWLjn0KO3HREw3M2h
KIe/73VQHrSB2hv0llIXv2110vspQYBYEF/Hm6EX8ffys/jjZlE5IBcQZUvx2YOc
YquBIbabVfBmX+ZfPBeKUMi9dni6fs/WGZbKqW4kjOtQVSCJ/gfiw3ki6UbyP/Lk
9kWToFSDxEr6ezuWSE4qPH73vJ4sqszo8sOzFAEOkjPhNvgqLR++KDSLLOnSCVhd
EuuL/yKwVjrZFD4BnnU9Y5YdyM/QSWOKciaxOYdkIurNwf9YCVBU6Ch6LlwUmLFW
X2lp5zlodyvuLaufEwv+noEPYWD5wLZAa6aOal/HWWemRmWhszRHkrH3aYiZ81Dl
4RWUpfhHQNZKP/YD1AIZ+1BHeoXLFkyU3xB7Z4YG9f2yc9aXddNvntknVRv9XN3K
31Y/pozICo3XV1/mrb7G0hc1o9LDPx0tdN1S4ohIPqdjl6TGg1A+BK1XuudHLVH/
HwNDHlChwXRGOSOmI/UT958jAuZ3Gd/8+MutxMttDz3zYrp/GY9TUVmjrQ+2n/aK
qiJWA4cM3AGi8edtDHTXHph+BMPO+ip28nDvOPe6D7sMfIvJ0gka/XVTolaRSvgG
LYW02pNKjxKGOPBB1aPt5lbjs6veoTAcyDhSbLfTIPz7h0wEs4mMGEcmB5UyCAYr
BJCNWlC8EVQbr/bF7RfBr1/l7G3f1adr3Y8ZlriMFoYG322ncczgLraQAHEOguey
GbS1uLIBGLWtYuelOx4NZZwcHhnpGBa9XE16ZPkalTPDleiGc4O2DKM1qawf4nGY
f/8IniY8seGpdk+MUldLJNZ8UIhVA+V3ocpGRRZAXf+JsUY5lfx/WzHsjaH8AArQ
A/RkGQqIjB0gkW8Ya9uln/7Rjizy4TYBAZF9m0/iU+5LohSnoLQL5+4JL7/3zYyC
T5PMLjbBnjWS+x2h7mFipLMIfuQBEXpauikuQNPqvPjiAjhxS5jcc8jjZTlJcKml
ddNXRkWtFSSBYA5LVIDezfeJmLfCEXG7zo253tJhNIzthCR6Wkgsfggtwumz5MZ5
g0jn+nxI8jKxcUUWKlETTfYJG6RRqea4IM8MAbn7dpeFxz82Mjo12+RFl87zMBX4
cl9z2pVblb3/fByQD4fN5dgUTyfeVG4x1ZRW/1OGSXmsNewsYJBkwm5g+yKuQudd
x8xwuNNq1K1MV/usBRaOIBzqtIuv7oE4P8mSSM9R+GUuXO1ULF1eUpDZ6Oipm8E9
BAK5E9snjg8WwZ2G50pBy+J5uZ7J6ETFT5rpFmBkRqQMAShPGYzH+aq28SrW3hEG
mcnBHrQ95p0P19xJ2ozz3KzrGqiuIU88IaYTPkJJq09HU0M4QtJCjrSWu6sKoFET
4q3Wl/TmlQzs6n6gmgSRxp2mdGz2nGNAczJuKuK9FXOH6FmP55a6/vZJN65/3fp0
toTovfmWL4wM6oRq6I2t7Zd21Hu29xx9eabdFyBJ8dBnOILwjjs85Am9NBt0U7hG
7Z2bF8JjLkrcCw5H1ZMx8rWsY3h/N6UZRZoAvCP9STrPTUaOB9B8XMDNC/AZZdZc
6W519ck7+zK9Gm5ARWtyl7ChH45RO3nPgiTqWJjz8zaedusYKlCMajsZpiWcr7RH
4yjspZDVPj76PbHESbQ19R5LkaGE5kev+rDhtQgIsGrZwAtHCcVAaDGTVKdpWJRl
6B8rUjYK9rMD4OJbTz11BYsWH9ieoPoxiWemyUxUCK0cBI1j6zbv+87ju9iS6XEW
XdIvvVEste8IOnC25FqD5NTRSwYJ0vmADvK3iRL/ybv7FIt06NbpeSMwD2AZvDfk
JElFR2rKGW0zuZQYocwfATNWhWH55wkT9wf361MjRZJq32RseLQptS9j+Suo2BcT
VbdZx3phcMOJ2r41U+sG3BfhcEAjYIacoFjW74krv6eokD2a4mYEcvvJqmGCLp52
l0+lzENT5cRnH0njMYnD3HTx1m7NfxZChzFlcYn6LLrgOOfxbCoR5rtfbFT10WRC
fwTIBJ7iBGiaNx6u+bhiLhMxPXZyVS1ksCC7rRfaRCHoFIS7JHgzADR+EvoHs8Ih
NLWAqyJQ1RVtYOOymcAV0ZRdyMqvuES1lMKzoqiPSHTQnwe3hTfxytBunCuFvv0s
TPtiBycu2Zv9RmfOgPDoyXUs/hD8T+zWlFU5CJizE1J6coWytIbzsERYdtEAfOOf
1ScZbdHatc78a9RdU5+Egc+4LyLh4g9lnNhbryTwVE6wOisCA7GQYBFhsNXUCYi1
2r48ncx5FUBGDLzHbEr5VjgDgPAHDol7q3J8jlRqbOryE9C3Oy3qaH52lMODaEwb
UBDZdvk0hgTwEQSvmZbP/nKvghmqB0vAomd//R2zUPeRrmPu8bK9DULtZjXi+IOU
OWh6FAZYSHgNbFz5xWntgm5y/75FCyZ3Xq+Q6wR6O+oC+XHeKvaHDd+j+cwwEmDa
a0b4Th1JvIEwZdMI5XdyrqDOMoicPIKczNv0nhJL0VOaLkMuJZpGpGfSz8RXXtm9
XGYhls0T30BH8JizkDmUGs9Uxq0JAlJd+Nf7DvH2HRLi1ZwHgzEGbSACmqM9E0Ez
iv3Bc0Jw78SYQcJ/a/7izCEweXsT4AxwehSKrUhJJtVuGvHPjjdcUqWQQ8LkOS31
WRl/LZynIhtT7Cb0oaQxZp2lxW6irdaFxlLUrtKosD76k/hvXbv2TzH3tVFyLgqb
no1qFuqhXu11Rl0C3p2omvvE0f1ZX55CDQ4kTM1oxUnF3OgEAkmC9XaqdLF6HRrY
tYj6QPLDSpGoPb9jMbsqLapkUaZxUAD/TSCV9fW9rMuQIQT/yrunJ1fDXIZuGly0
x9oIMpgrHLMmkXptli05w1qnECPEYfNb/kqIW7q7N0ewTiF5f+1BEcKZnly/Ocm6
chrh9hgnWJZwUtzFmpfTgrNJXvDrleK6VTLyrxd50O24IAq3mDquJ2T7s3iGr67X
isi4XZmCQOhm5ZxG4KXidNBqX0vFveDEXN38IKr3oOaZo6aqJEJrQubi6UmyFB2S
6c87epsuIxm3Ekoezg/VNk/RtjtcnrhC3uFeUfkRYGTMLtC8ysNnHnWXXBA4wl4j
+ceWQllnOvEFFeAQeip0vl6pSQSTO2N/XkjP+nUm916H0n4fQa24vpEbJMkiGUHz
txvV0HlSaHbYBlwN7/NKuj3/nAU7PFnHjbYkj665/5Ef5iM4D984NnFysyqV+2t+
jDer+A8ZHSfUEQIPWKVzThmM37VlEb7H8NivhfVFFwXkXcJOVVik9p7qXEpDbjQZ
x17SFGYHxNI4rGqo1cZurxL0C25ROKaLiqp52rGX7Z8Fqp3yhQ+sn+9LnHhsCbg+
ziMQ58zByD2ZytWY0SYjbNQGHH3VQDMt0rTv06uspyikUWul5EoKWvNqzS6z7MIA
BTfHWT8xNlr+NCcBzJ5FvuX/uHt1k4BcFKGZMdG1K1R0vtykrPga+llq6g7hAwjz
OFzolNlke5pB6X6vo/vHpyiFSFEvyNANYuv5ZLIsVZGzFFap/6TUTN2Xcjenk8IE
Sxwzz1eClWShjuCabjhrUkxu9MsvP3nX2rFO5sZEI4J67DG06CrtgQecTSPCx/UD
4AaK3LPsEOPn2yrYCA8iV/NAxVZHgOAIX0SyZEQkzGpnZJwHzvImVL2ObvyA/a7X
hIIDUNc0XorLf7PCf60gIKidok6WCbd4o1Ka+AZjr4pB7l3QUg4rXp7AlJVc7a6p
Thy14nkG95jGpaSSSVmy1Y+nyW/DphfdMXkCYUWmUOsuXpxwIGVJYT01eVZTsJhA
U5BERxeOE9eoFILm0MloxNlrZNBQLwZ/DJG1RfBQtkMMmADuxbGAy24h/tHADcLw
LWrQU0SNlGmbmhLaBROaOPp8BW2O/KPEWzKBxGHYgq9Q2NRC9EmpwfxhnXsmmayR
tm7YEuzqGMy9XaAKRD+aSjLTFC+XbIrP+TjGexYgv6YtbBZEWpVB0tojwTA5NNxz
vqJ/73XRmFhQZqpMexQQBoWzXbALyQedp5QRQzNatCXaulPkqtEdENQRxbYRt7lA
FVmcdS551ASqdJllb8UUhRwpdJDiGEqveyO4l1/k3UkkwVZ1IUOJEOyIbcjnWkmY
IdQNFwRYV+z5bXvQcdNysdYntHi49Vci8J3Oo1YsfM2XrFi3Qt1xHMSGhhEC4uZ+
gEn8SCyCGafttIX/s25SA3w4uGdbCl8A5kYVXms+muLSxXAt8pKoBXLi9I1FbY6J
QLSKOeT1j0oyocSSL+BR1M4lbYjd97FtUTHn+vOsUV2mFVqOaRsFq3vcaXCcpiIE
4m2PWPUiuvqpHe8D4cRbyZMEj2gLszXNu/g/LOUvdkq/sVNYyP16QrWiTPEfX9Fh
/tiMd4QEhNHPANYUdsnK4EPNa6Hc1K4FrfIkjqn1+fRMJX2n2JGYSaJI4kr/Kt4J
aple1keM12So/v7SaNGSci5g4hpR2q66id5bfT6rZW0PJ5b6eAtQO2Gs0VF0PIn9
5gKKLcAtPOxkhc9aOSpkUeEBW0704tID9X9leYEhAG/T7xI7cU0DytUp2RfIDMSo
0bcOfLc5oRFccDoLKUHm6Kuz4FNeST629skCi+DirjmzdpCxZKCF5rzMaLxV6DuJ
AX9A38PCCui90aQ85v3G9gXE7D7R8JLlLmIaZn+VgUc3NLqEsPBuLBh/wLaOMnYf
ABrsKzK0NjuIabVSlhtXgvqSuI3eRWMi/xbiLezWI5tJvM4UHHXxiBHOh8ARhcrP
j8ngZO5a2z+6bkNnoXiYzOpm27rAyQHUoqpfII55reR8ihXEhX5BiDdWGGGI1HGZ
TtBVppekIeAfPQwkPAiwOPYPSkzeVBJ5jP3T85CHmlfvw/wEu0zd7IBjnRKoHiSu
TLB/Cm3yWkIEFh2/wMh/8FE9sCaOx9peZVMjghfBZ9zN7/Th60mYy1g1qmDInFlH
yk3d4kukoQFiB1bk06iHcZ7MCeSQXca/5mhGNSsa5O4/UNeOWQz41fqyi5o+0hPX
osD02KYhgyk9yEg7sr9sK4+IhhxxLRjf1S4/qhl0NYGLpW1WtzudfKs4iPuX8k6L
+NhhFdcBnoF1ZeehCXutbQOQUSMC2KgUujZSy+EdNU4ck2pzBgLOY/q7Ojg7Lhzj
ayV0APbSk5rIjelXpnnjb7Q+BRVqxmklUVKrTTR6tAlznDnRoBq7YR0/bFa2rPKP
0jkNTP3Bx6cMdaQGHVFTTLfNCdMvILFXd6r0Haa2QRtnL1BKXX08Qiw/n81CIKst
BUgyDlVnims4iIRMOMnZ5NXVMeyJpvPYkbRIpoH2oSYDHEmVvQVxqfZX0h0jHBNA
oHb3U9FH9vwCUf7xWjRgKDD/gdi6mluYX5LWi5t2f8IUujRjkFSCo+RyAQo2MV5L
Qafj/GeNDu4QFfsrFcVjJnCrmxGXmmJmy5XnNPSS0lJbHlNaGX6Szv4nSoNJCQEF
4uAd74+eE5US9oDVpnD3/33fyjZH5OrOeXFxa28cYdtQon4iQD2JJcdYHWxaaLpL
dYcnPUEXYqESJVFxImsGYXbtS1LmaZ51Vmwl+vPLPvToIXPQQzb1hQV3y/2WgGGX
n31Pi2PZNDBwTAtrIV0Wb3ZJKykKmvpGph6yh6zjqH+qwb4HAuNM04fsaAwJSDKq
HA+8bYxIaIcFVeKpBuic+2auxd6UJaVXHPEuvPlQ0lsUxxnvPGdn+80Yohi+nP9t
0WXKLM8msHwmytLz4aa51QgxBKcngxBdMAYuN1ojhWMpyi0gOPkkBhjql4VRped/
pzRDq+B0DDjJv4YsAYgyNFPt2YpTET3YTQGEdTfWq0gjYUzh1smL1N/P3xVIu0QY
mbti507jSgNeTSYDzDwM3OGyhgTJWVUJDiCIK7rOFIfzn+lWDaqwPxkAl3yQ5hrc
9+U07RAEmLDCjubDbMxRym4VhL6vbK7uKlIJMYn8rRHv4I2i1Ux5XNgoMgUAqs6C
XDrUdBcQmLCluVmi1CLnUu9NTkAD7vfzlN5UQ6YOW/s42zSnE+f81l9MX6RCPkhf
7DNOsTIDh5z4s8HgnflwgoTHL1ukClc7OaNQdTbE37x3yXYmxBQHBPlck3usOjfU
Bt8OwnquOzIfZ6457DPgQ5LlDxl5pQAzD+R3OcLEuURDDZETh4+07A4zt+N0Vx2W
OOYotDdahmn4nZmR8XejecBf/76IPUJz1p81Rs8BbgS+pj8vA+N+qnCDg+A2TPvs
lx6bbTh1v8tMsweFoMpTzQwlej1pz28NmqvDlGl1cL2cSgb6R54wkkMDOC7J+YKN
oLs1GsMXmgMWJGnYS0YgVkdk9xaH0ReGDh5fq6WI0yMVjQ2OqxajKxoFB+DtCEKt
ifH9dDz/3q2da6Rf5lmFLeG671B9dwd4Z7/XhVtbgLQwnVLDlTxS5OdkRNiZL0ZE
MB0KEObZyJDQjPoyQaINtFA9r5HNFdjkGauMrN948pEMInaN9FBjIeYy16XOXKcm
POfyQnh5T7n+6ZE8mns/tsbT54jKU7ZRMxdr4zabp96Rqs8DHoBtDjsR2ekAJe9b
MYS02tmVfJazW3DugO9DHwQdX3pO6tYLHG2s5YFpnkw3C0qG1qDXgUvjY9qIZIo9
hPeTHFsu0MivYwU5zoQ2QKw21mGqBnuoNg4RDi+RsJ4C+aIBviQFemR7ADdsF01M
UZ4lt06VKsr4n2h5kWYep0yvPqf83at+PIm+DcsINQ3bVBDcwyH3E9bBSiwsdxNS
qSQvTwCBmq3nP5CYbUma1ucsvHuBNufvPTB4JAKOxQVI8sahtEKF0yUuXWdifaJu
CeYCO46yvInX2xNLKBBm/mywd0YLCND295bHM8gu1X9/bledU9F5tjUzGE/km2km
KTSQ8ZOjphoHyMVVP3RklohQGoPTVzZkziLedMRp17EDywIpP4CdfiZT1/8huZFd
cyonuqL/0A0SLkYHEniW2h5n8j8FRcPH9OTIsv6urlgGVus0uXucL/gVRxOWNHkl
2KCQYjVEL2pitZLyv8SdwI6HAItVlgNahnfNLR4vYALGRB8N0DNW5xVs6P68QweW
EeaZoiCgiQvrOMrPsb8PTW1SSefjrd8pNsuUa0dkbz/sCsfzRmG+f+IRdMu/vEg4
8eEysnToFS9eY5kQUla9EOneM091KCGsIB5I/EKQMlS+9bMqkYfL3ZhNimJmyRXG
bmRSpLbHSffYY12IxT69SO5jLF0yo+vIenn5vQR38b+fxgs+VqCg0wwxfXjY5CxH
Np1A1w7kYAj0aUIIAE+4RG+clUW/9BezJQ+Jzjpb0pw9a/+IjtGDHXlFiPJtEET3
uHiq7cXq1Q8lHFVM7GOvJNja5VwLu3HCuS7N1zdbdn3njAEFtfAHVOa3//QaX0DI
kontjgRNJOlvVRtyvY3TlXRGScteLYc/Oes+/0GCe1tQxKC4HRx7qPlgOkmRUg8r
p1INoSQSA1rcyRbcg7aAT1+nzBytSm0Km2BqYapIFu7onsKE3m9GxikAXRfEUSb5
j7dtx4Af/G+f6XWC8GBXWqz85Rp0tWzjXMjoS5Bv+487QS+4KcH0YUJX/XIeBXzF
L+8uTytEzoAVNB1TgM103fR17Vv17yyeliA2jJ7gJmr621od02tquLro9M/T5vHZ
ZXDs+PtIGHsRVdkxLAPO7JAxuu2pGUgWXtHJU2BSJXIkHd7dWCFOVwyslWnsFs5K
cd5scH87nAONfc5toQLqvn6+pEshh0LGFz+Znf3u4DNq/eivyVegoSLIyM5SVOAP
nP0yxTYD97qFW+8LEGrrSdnvvj2C20nO5jcKo8C5kP+G6/emsdTpEgTrJwgxAogX
FR50LGgxmcZpTksyhCZzKU27QpGiI/CwzrFbtuyvoPvjeBtsepP5gAXJey/Z+lad
/5OETB0qg+fbTnXqvM4nXp1DBJ7v8RScbWkoVkoacOJRcpp6HRmrTBlGt6DzrVzi
y00m5T5WAC4c38c9vsawf4jYjIhCa+Z95dIV0IlF92WK1S/AaxHJK00ckKBmN3QK
7nO3k0Vud6tpZBKmoFcolayGsE9U8jBJQWEnJp2KaCFe6BoEHimR1x4aYncfdYMR
jlXcI0fAzzjrwrgMPoTQxajSyYEPFT/wTLk67IkkAEh6nhCjlcHBBVXpAIENOR1L
k0smStfE5fE84VNkb6Mkr9CXhHNlYOHwOkkY109r1ulJErKg5yEy1DbkugJiYoX2
xP/O5XBGMiVOGQAsv3sXY2O2ITyTUDPPH7whHflkanbQnwLr3vL6vSQ2GmjSTHZS
dHxfKa8qYzRqktsB/lQtizRoIDMwvNQAaOouhb558G3SSJnPUd4qmBGzP3A4gZq3
PesDZ7scmtfubBmw6DKbH01iLPLIxI1Q0dpKzY/X4+jOh4QW6l4oLSKQkKM+8Fh5
pW99cRe+R5hkcO1JBrL7UZGi/7SE1ycgCv+PAWteYqm+7dV1bFxec8OpuxuaIgfp
jaIppqUbWMkxZgRIv+D+5ybPNRgWPAfmDyxyuHNXL/6aZUVW2w5SbtGTI9s5Buk6
t1H7/tAZmN3PYzOBnzqEUzjgQI68bZEJ13RTXjQrEIRdXk+YvaFaM1uxqii2brua
Erae/31hYZpp3ccPuRCBTPTrZWYN1hc3d7gbh1PPPqVgsaS1Qd8FZbg6luwiKxZ2
W2nfzSuyqQ3HqAXAakEYl5u7hzKedEvBt7eVdwxFVNxC2Cy8JUa5ztEe81qtTLVZ
muTEi4JGkRqSlkwp8CxJa4GkmOMutCGmOYKed9UdJZ1gXaddtWYHHSbMgB5ls2wZ
QTgiAWe/6QvqeniqAb9ru7vg3f0F+rNsT3N11IqzSKaI8BAjOmkcManV7xlE30mg
g5CAd7n4zmErFBOwbJhmJclY84aJHXwQh3KoHcdWRstD+796POj8RH0ct1UmiUBY
+4gJyBuhbUE4aJumhijfMz6OuKMXEriSQnFMAkj90q4ALet1GHTH8rEAPm4OTbml
rw/zjFjIEeGVshcEczNSl+vUwNM+6R/eqs6NmSd0gAdY7jBgFN3RD4yVss7gr9a1
1VXWMjcudUyBGozvHOdZzbjKJFZZCPt22+zjQfPt/3qHeXK6wDcy06ahm6XoBZw6
l1NSGYQHeD+kAR3/YHjbpDNi/w4iaUkh0mrbNFmbNpF/AcjpBm5CkJRHtPZ4MRoc
tLK5sxLeC4lFnDXSmrEWYwJgdzGByS8gB4mz9vBbyroEIx/ZsgRjsjclqvRKE7lY
FXIAbDZcY/P3WWNyI1BlKNU3x58tEjixW64DoaytHSNlPjMikxTzkNlt8Q96J5Us
kgrgKOXpcjnTi8XT9RmK3CioLoLUiw8eh7D8fDO7l619dMUS1Abynil9J0UuNP+S
GlgLrQh+Fk6yg6gghjCMrgpL25LKnazJZgDUkiv/7bqfA191aNryMvkLBnbB0K6a
aM8g8Yk+GyA/4+c3YJTz61laoFbo1mvntkG5CtfQ4V/xJNyxbHsK7f4zDamn6t+C
pB3AAjfchxAKN2PlJLkGnaY4RrxqBBlV2xLcXwDEqobpQXbx0SWdl7qqecpBQ86s
oj7j41RYbZbwu9ifI8sWohIWkykDALV5lfDVOff3nBOflylz6IPqs7FoXdBgw5qo
dKLfsuRUh48Iemw99AAbULg3+yNDZAFR7NLRfvEwM74/2wQaErFJKWbIJE+sR0EK
gTpcyOBz4+GDwoSQHxDXlfsASSZTuh2jEbgQIbaGOdtWZx7PXctpv3bh2N3MLfGI
P3/lz9nwsa4uKUY6bMBmhCAH+ZH5ApXz6QGJpzh9boKGz6yoALEnciMNJxyRM31n
d1gYsuWzvVkklzKFzipU4G2TYRSjqfH8Kz2NaNdEbfcsOPDFJheVxf32XSKvGo+i
JLeekjbdr6wYt7QHjRsntmmSa9vWGJtJ3QIl8iosqDzJgE5I06yFSDNtwPkYmCvy
/iadDJHvhogIIMgjTtTD/hSZfuoNc9C8R3fevDawo3NZCLXSVW4rN0Aj1hXtot/q
YcGUm4U6buSDpq9yKAtIcSb8xGoV+hrrmqxwp9E/GR0YuGM6KnSCzMNchmoM0AuK
mirIiuVRFth/uo9vN0f3DphDYUf50JSxeglR4nQeIdfMNwARM7a/pV3uat5rAFFL
kSmihE11VESwRSR1qd397/d/j5cRGOiY1QSHpm+j+bIA6GT8fH+yl0TTawsU55jj
IiRWfopc+HQFKaWbe352DfTnO7VENHImW8wLAY8tBnLpOcLEdbVi/6aLc0FHIv6x
/y1G4APKXOLB8PE0SWsC1Qk3uADXGPg394EHm3n3CJj+0nfqn+NB/hw2gvoASeli
ilncqDKL8zbhtcQeAm/XlG926RiWRtF6fKMmMweW//7fre2/yr7o+prY9DbfIIiu
PgULzLFrnf43TzB0PSGPdPpS3YSirPji0AusQ5Z8dnVSw+YnFrqmRXwD05Nz1+oV
9apTc4j5NPBnrWqxW1gGSi8apgn9cufeiuk3neZ7D6+/kR+jVxIvGrC+SHRNAD4Z
oCidccC6mTucz6hui1uf1HrfOycv81d1RHFBOdDA/cvEEhb9gzZXf+8yK2kjNaRz
7JE0wKMmFnT9w6OkotWyYQ1Ad9sR+Dmhz8GsbcSAT0PQ7zWb/+h/MrYkuFREBRCd
2WBqZZV3OPJDGcNVh5S9YqNUokzULz6zLhfjeVBlZu3il3EdeJEhSzwgupeyy0hf
WxceBsl41za+QzAkJ1JbgZUQE7aVavTi6eQInmYU5xJyAIOHliJP6han5iHjWOEh
bM1VeSBfcvOFdCQ3hNEd+AvCeopnvq902bXvEL8DIImvCWEz46lpNnuKbDIGyCYg
Wnn1ctyVKWwa3zQBjA9tIiriUnZUxfOodq9N1Pv93Ov9IOQALLdotoxv+u4ejgRP
a0RQhRNEOmAp7Xx//QGr5yY2NGFsu4HPI+M0+tzrzcjW8tJroGv+I7r59AztRflk
Z6DQb7ZP6OXc7Yk3RoXhmBk4LKgQpYQdeV0h2ZveJ0p4dV8n07Xs5tM5Td1Uw3Rh
nsJ7X/D20TSAkcLSOF1dhmeTm5Z9KwiFOIrp+OyzCtmg9IokIuiC1ad6cnpYe1pX
q5e7kSTiSGygux5wsJBJXdxFbo49rAw34TFAlppmDyDqzzEJmxPjy0y0LnNw1sKm
5RjwuMsF8kk1Qu2cR7yPUEVyeDKOKBFr1BULKz89q+wvi38ef1u10Zk/mcG66C0B
+e91wP1RkZ4BVcnsetSacSYLe8xRL1RRg8FOMJsAd0u41vr6HziDo7NFwuX3ax9e
Vf+ovQbdEYuDn3h/gopZKNMPSn+hcwIZf+Oa4J40TNGCPe1558Li1/qs2/zTVnKF
6+nW95g+3wUSUGklDkNh1CZE7EA/rxIx9GlLpRWS4Tp9LG2dnOmg+LfsKxVXiJm4
q9nw2euCV3+EYnwyTncZxmY7CWdF9pUOp2yiXcwdhC9F0p5VD9Ybj7lSAgTt10ko
2pq7tCBwuyDQo9ypvHc7igSiz2V9pkX2QhcW4kSKWyk/dF8snBaBBMt2eVsv+do5
sn3nrTnQJ8lmJpjFyg/R4k6P271aezrR/BeyIcs2h/jXFzbOhe2/9wolIbHp31qR
wnwsasFMQFuvC9Ni7fpSPtDyrgdLJyABMjNjdVkBeosnglm65kyrz5RCcVXeW0zo
V+X0Phg21/U7Wym/7n6iDkiQ5i/PcM46l7yPaZqk3Akr7vSsGGMaZmdhZBqexo4Y
DequXNtWfp7ELbUABwVQGyq9B1PMIxs7I1+Kc7QmEtDiEzcxiegfFdsOFEwatUcx
JwYC0eUUb25aEZ5Njq2bIK7cBktNCJh4YKymRC28xvEifBuONro+dwwnXCNznKa5
6ao+HLU2/ascUnNCeamdawYRlZDUBdfz/ZSAjtK+nmeHO4MEk1t44xUfsGFBi425
o513ZUbouQ+ecB69yZiEXNmXF6I5BgbjDmYiMP5TbW3hy8SwT76cRvJuocRtgBc4
QsephtOGFq+UIWA2aTo0/l7z84pGUhVAunpbIHebrV0/WvCqHXNHpVdfXaN0X2qI
WocDWQSL5JHztmmiHuap81Xs0ldho1GzWmmFkr1fZODR3n5IiJhVJDDNTrLoCaMt
LjcLxzjt11tQbcHZ7sgWvGiZzVe9suqXwrUZmzgNd9ThZxazaj/pAhey/uy89S3N
ysS96/ibdibgph+4wfDyU6vrQt67//XtBZo5movtMKNt3M8MPk1PC+9REKEl6p6l
RbKtSL3/7Q3h4qRv1NqOcGNx5RhqErotqLVZ/tES4brZCmiVF5vyJRYJzV+wdJb/
9uHVO/XLMUV601gFPiz0t/X5HYydXdz/FULaujIRbNHjBD73sVynAhYDTSaMisay
rapHPpVDjOllFmsbq3Pu5qc2DSV98bjsKCKw2S5N6PRaUfwf6uv6dzInaBDd9Lo9
/G77tKGjgZmtia6hgwNU6wunQG9wuCpXZwyYa2LVqtC3DgeHFt7fXQQl2G0v3hlS
N3U6Dx9kfdRQ8K5gx9YsavuYcMlw+9gki+CoVzjaYkNEXlNFn+afe3JCpXU2kNWu
KG4wuLjwYdjyxcSSvxJ5u3IgsgcInhK6n2gdtyj53Zb0ck1N3OHDRgju6T4dEIkI
TB+pMSwATDzHyt+GAYYbNkQ8DgQUe6yFLS/eHAIh9w/nweEQqayP5BgOp/+WUL3t
6EQqtPxShvP9cJ+dDXJcbnlXw1gkBhk/qMEv03M+/wx05sULJvCYLXNx/dRBcSWb
/JvFs6+Lx5+POrDSja0Z7z9e3shvL5VTpg7D/juMFAX5Vf/TzXCz/QAzFnKnvZ1Q
IgIlYSIDYEz6MQTjYjpaOiNGbX6nATjQ1RA0JqelkfdgfNXWPKJbMEj/J2JLM+GC
DG+tba/jFhA7SDOuYQmbto8gn8/bucDM5RMbvPw1V+73MjJW89Kv5ukPwWYQgD3W
JhK45Wgt7MEqXym9rQRmCGXRQCmG3ZFCg5tdC19MCkP6LFW0B9heCprhOWWxoyu8
FRM/edCAh9gmaajnxhCXTkIqgI/sqNozPaSsbRdqN6QEvCCyhJ0ExEWVBF12nVzB
xXxrryyXrvGHvp7yoxhJmB0BIIJQyjhEohsKtjRu+eNjs2bihKe0h0Xa8mYHRcNW
L192/BuMY2+0Nc58H/fMyskkvxPuA2CMPHsedPrpfB5wGQc72vUO0/eFLqqWuYEz
1KHJ6W9rPCaZdYD1m+Z7d0WU2FC2eHh1XgTh6lO0VIXW8eEiZNGkrko6u6W3d86L
LjO24jbKv9BZDzfxE4jkNm/1k81rS+o4T4kSeZnK2YoAyTxRTa/MDeAuRWXlSjht
Q52QDhfxWV1xGGfC8CNUy15HzdePzeIQm/n6KgYxt6bsI1u6nHYa/SRbPUHzAO71
Jso2ZFviCZglEiP50tkkjVSfOwBA7QFXYRuYDfl+i1eHhXXfq+lbIUIkOLnlB2aP
PCqcHzyYfrT+i+DOB2gPSGDZxLkbSY167yr6WKXweuxHeyOTuANJKbemsUaHsR+g
sMIkQmWhsIz08CYMdn6ubr1vWY+rwZl9CfWK9gc/niaFu1T+H0nv+GKweCiUsPMv
reCHebhe9VvuXqx6zZSpecg98qZZibcVxSuX9UkUQSXYWMVB0lvkkFjjkCaumrEu
6wIv4JwKBOCKdCkklIB1p1UAxFa0HNiHP7qxXZJ4hh1bnNj0LeWrDPwdcdJ74SvK
pYnkL/yErmo2KP46fhNUd9A8SJmflgoWUbd1OfpMfCsC1jetwZXirhsZ67p5b/py
fLsz8OG7wfKwZZ9lodxifBao3E4lFEB+uyeCv3K9FXym4bay2qB6k1x7tcXsl29G
ndQGMNvRXeVkOv2sbAwuThhkceL5hVcHgDWWiAKvMttu++yF+DIzvreUW0xoo7xZ
+oYBbDlmS+jIldOrQxLlDE8Rd3JkIATIhZJ6bjAWu/B1m5qnNuoibtIgGxM1Z+V9
F+xBW8hZVrtmuvQ/IFTFJFmd0HSCldMGv0LupGZngtne9ehmo+5ld6oD3hrwo5O/
qy46K+KNzTmnLgxlBwOPqpGczs+cU1S9Qcd00HooxWbj4CwNihFRPklYk64VopYj
/t1xh6b1Un3nreIGWAzN9o6t0yA8AzAXthkMrQXvDD1/z79dftHljXL5jmMkiJeI
T870p8hRyFHCp5z3PuM9Q2o8aDSP+E5v14VxpJz0Za4BKbaf2Zj5f7zPiYKa9JVN
pY3v2zPYIBA4wy0smrDxBMv4vu2Qr1VYdeFUT60Yi1OXtcJTnssSvjPRIkt1gK6c
ukUWJEjLdG5HGf/3ei6UVuEHYDSpj7tCC7VEVcl21cz7p/pM8WoSEXUhnVsQtDHl
D8UsqbFGS14CYbkSMY29k29uIh90URI9WhzKPQm4hTshWyVKf3Nz2X7SBwWU17El
xRR64K4wP/pkdVx/mDCq6lwWWCNW98EUqM7ol+L+CV99D4dSg/eOoNa6XImd6DYl
n/oTW1IC006U/NBevEJoEAlXaO7/xMqrbNrJJAM5eZcCIhGrvQ1MvNHBrp6aMF+1
amUBbFVid2Tatbl0MzI8JdC1KIj7S7gp09xx4hhd6LcmwtK4En297muOZvDveJyJ
tpFwQsTlYNGFfraUD+aT8iCRLIMNXG9/dxDwTtqUXYmGuch4ED9o+Q+oZk6DkGw5
WEmyqDFy7sKLy3jDUVwFpQq/ZOiyDl8geAAcbsHugJ4RjLHymugn+fLw+rb/KC9K
mxCu5eaRsJYJtvCrzWi/0a9SOkN4uzoVTXkEzgyPO4iEgAP2zx4r77RyzaSmlB73
eOh3/JQbFCuzXXc6MePa4LUhgs+VOMRfiMHs6ayNyjF7kkeoxDZOLGIVU8qcBKmN
/YvAR5hCYBPksxxukwn1qHwK510Tu9IlSp8ggkLDUDJYhMBp6ugz6GuNxZBnnhRi
LD0mSLdo/13LTu/dQTNCBLe1d0iobM1tlNDcGon+yiNF0EqUk7vu0/ERdG6/Jmib
e028mF5D7tY7xKjklr9Im86pp4dkf/54wZV3FA3l4ZX8il9NOkrR/NbZkV1Lt38N
lvIeor/4DLdyoMPf2DMqWfaa0CE2XxyGx4xe5rPjZidgYPILBkO4JoIyjv+K1ZvC
dp8nJWGQvrzA71p2fCfQcyli08LEhBtIdg5sgKaAU4aGWeSUi6wIQN2EVwNtZ68o
1WQCdbHoHXydBPOKYuxLHqlZuCyg7mPpJqMlKD9k6r7svc2e3x8r9uR/8u8VE2YL
MZHf6uzl46cpBHQCzEtrYCbpSMJxbePAxiCw+ccy/6fR/MeelHXdIRIFPD5nsxxa
7wKicZWB5uNO+wwhC82AkDqDzdXuUc9tGyDow0WD6pr6TjZldkPbeOJJ5Cg2N3ar
PlzVVHK8yZ6ifc6WjZXWYtfaQXj/Ex3tiymc1HB9SeHRR3CXMLBMeo4TKhX8vSap
4Bhve0WI1kEwEHMjlgedKXSLPNfkUa3qPPKR1hArJCod333skzYg2L9j/fjM/c5q
40DnVr+3LCw05EOopSpqIF9bHSN/a9vQYSShcSs2Vt+wHZZg2mPS1MKP6a7XRZPG
UMdYiV7Kr3rTXKZQvIHUc0BPuA88I0T1rDVY9XkDsCAiBTIEGsJV5RpUhxDiZ9ix
5sWDC0qSgu23egj8PUR9Xt501vPJFa1XkzkxF21dIipvvNOIpkGKhODZHvyPkDEP
ZltBGa3wTyuLc/mwtMYZSdmscHgjE8EdWJGueOjiicNNPMU64lDKffCE3QBI6sAv
i9qwGSsfXYb9S9R3o1jsdlJIPfhKdIRnDcZTws38xdQAXX2+PyKGWp/0ClVg8IU3
5D8P8DJi6mMNZT4Y4dvdJ3HeV6EvpIBtxL4SWS2czOQvL1sKje5QWhzswTCCOShu
CoWEZKOvtSqbjkQGNs8MLfxEzGlb1Flp1ITsgQH6OONf/7HikUrmu1uuboG4qPQY
chpcyX64OUmx5nudtQyM1EJAivcfIJh+OcAG4bOOB2eOyKWPmvmS2uJ3jLx3uzrX
2IdUGcp0TgVAky1+36mDiJtWMW6Hdw+phyWmkBmC3yZ0o0FG1J6soHXGtvKaleUh
Lf0UIWE9sjt6trlEnDc6lu48UnWxroNUU/54OPb9DLjCmgL8n6RM2N2DGXl8hklW
EsN5riu2HLubLpGW6EWHrViSfPRFe8VibLa6VDGCZdIIpHvGZAW5FqUGcwDHmKYD
oLhckIGZkLDjGCAazudn8JatzIBMbC6tBoSqFJaVZJfobPO+f5yJl2baNLhRCTW9
qLdpEugGwP4U2shxPK9B4Ly7kkggi2hFjJbi68cGxvj83YKDQbgf+kq/qhWW6zig
rdI05UhHC08cGcuUTIYj0psI6s75tsQDeTT14QiSOuaaYtcb5IAidEKRP/Rh/3MO
/xsJsG/kxhc70PMlFqAXvs5RF/HBGKUBO5B8yLO2bFc4XQu39s5e8Ycdd1ZaeCiK
HJWOH/fMSZmn9kcUJBweoMiC+ibPFEvgluXrA13/xX9k/aVN5qUnrRaWJQtUyTH7
3IrN2CanvT+aQuiz5Kt9X03n3xd5iwVzYYVThAsGkwEYROa5I+Tm4aLKtB7DycVl
odCNANK9OOevTklpF32arqH149Ji+l7BhWBZEyfxjYgb4En5C33pNg5YaTt77ZvY
VWq9mqomiViaHDwDFOEQEgPj9X5fxxXNqFjRYJYsj2yCADwBcfZKFFk9Sdp+fukm
5uDqtccawB44XbFt1ryIF2uJu3vegJeGlsK/gx3gsBuQpqgF4AFER2JQpNRDLP/z
gBHudPd6NZUBLIzedovm0PSxoxI81LSTSyXZv4azw8/yOvG4cDH9d+RYLNb08HiK
NpGfklTMnvaIo7s9LVeox9rp6SKD69UxbPYKBmxG+7BUY+Qg914+P395zAB8WYZl
Rix3NEiLl3CEhtsO+II6rQ+S/LOGt2uRaogTmgjaIrzgrV6bvD0IX2G7dXURU5c5
j+UX/6WOkgHVO1cLQMFBYCgauRsuo+13ZvSDgqjJobTzdnI4RNbDL0gkwhSo0R0Q
o+bZE/I7gnnnD4I9DuYWhYzUoSKKX6B0y56JKxMR++sQuT2+Y7NEXfnJx0QNrgfp
nwLDnjT9uM6O7BMLmuQoPDwRHdm9Iwa6hedu5DAPQG7s5CxZQVk8zGZUV42jvkZT
jsmbnWbclk2jxwgwiaBLnHMzsLfh35rSPbCddaRxPvEzx12VaRgeSIslJq1E57c5
BqPC+FN1IPkW7wPvgBob2PltqGt7Luk0OLRhcBchoMFPRyG15cYQVbJM1Bx1RcCK
nqQAYK4VYjXAbgAEPZHP3fMlVdWE+13jcqOuyH1RS7XpMfVAAPXwwfwVtg9dKQ4h
1SNfUwXjr8X0vlBQqDjnFxIs3osG1OKup7+Qve6F3S1VCqcr7uFY4FoF516h+dAL
rtFk4ql4fHr09FT+5E3lDAGGWIdG7cGaVoaxSEA8iUblK3neTpHdtQpBkhbyR/rG
e/xuno5NSW3B6Z8GgwMse6M78fp0M9nMfJxSFfalovoqvOzr2hMstUHjFm38ARop
fYIRsv3mBm+lM7qDJBDxx7jTGcNzSoNP4zqYBwtseTaqF2hCDH6I9nTimOQy+UUE
dGr+0LKaXsVaJPkouro3bqs7QbIublO1VqLBR6S9CP8+UJS+/rnlsAmbmQISP0Mo
uGKO8qnuJO7chN2CGdnDL2S+yaADFacT5Pi9Yh5ww2pgszgHVn5BZEsr2GDZjSlf
DGJlQG/ionUVmvntJ5Da7VKMSifdsJc5nUa4j4cQ6EWkFQ/2Cbhf4w7ewvV3x7lk
ORKnsQ9OXvAnyo5FzKK0k8TBq8QkrDXPjaduFzSZOEYeJlMC2BuozwEs+KIbq9JE
zgR6RVJGlQs20KAONdC2SNwWvtxyqpOUofktbZyxrl10h+GTvsfnolZdvzNW5Jn1
eu42XJqqwC5XU3mG94bYK4VQKzY4jUx7bSnEWugu8BagQ17ymvvaAargeC3Mz8VN
6JENkZX9Z78PR4J30odOsPOKBWL/L0s3g9A1hFi/VptfW14/916zZ00gFt4Iy7vr
q84rvHzQXVUc+7z+gb2kjimZwuB2jaRBpjc78AF2iWlHaGGXBuKJV9EKABVKRIef
0oPtEGbpmTKWezzYgiNdBkVa9JKhFxFubqciWabfbeQD8wdPUosj92O2psNwGv8c
4brCzazxc5esU0yGG0voTwbwGePkmcNIumT56ffQAZWjygeb6qFPV8aHNW2bPPv+
CI8ZS1txrZkqoT8xQTcci7r9Pj06x3/40cbUC5iLU9gAIjmurIAHLQkGgVu81Ugk
oKUuJ72HfTlZrcFbMmjqurIvR5H0Z62motjDvYUSGtyNEkDrtZ3VypJUXMy4DGi4
q+r20kBUopF02Y59R4+KVqkXNzN++pFBuNM9McugtgcNmJgbCuHn2NQHXdTmKtlS
e+c/3LOMUqWsBt1zIKa1Tvb+arHod4HlNtr2Jb3AWxPqRm5/BZa9mVwBxPEnScQt
EhW5FEQB0jjNZeDzAbnA547fmw8XX2h64rGVylVWPiHaAJXiFij1njlt8Hq8Xglc
RSUSYfv0pplF8iDBZL9IMT6tcRDtXQK5UTX13VWvQ164Bp7JAM3VJyG7TQeZFREv
nmHATU5aTeCnWjdHsv1UwMJLAbzCeIDyEmb5gDb27dVQFJMXXhywj45rpNO2/cXq
QFABvrThiEsp/ja3lPr9W+TR4SbnU4O9j7x9NyT1ZwavQmJBHNoYNULFBoHTVvPp
JrnYEogQrHeoxkfQze6R7VBa7OO/eBr9ZZD0ptVAjPxed9xnbUXNzTfG3ELTs2K+
GIDbcKi0Nj80z1L73enXImld50pwv4kZZzB06kc9foyhzksxY+pyW32eGyaqQmr9
lKDrt4HNxO2+xgIRDGxYbCB8dMibfC6vRcsmbk3F+iaF7sGD2baLAsBisJQ1vXCR
afKICblyS1ll4kYTSxD1KMVkSruJMq7gQvOIA5sUCCIbZpfnaZrgaqUD5bIbnjVS
gSr89BPYY1bA1W+uE1IU9nXLY9FGsE2hra82x+5OVGRQZhrs+vxecnGuXyZBBPL4
WASka8k111UKuIgXYkTGfE0NmFTftiqlnJ8n+cDXQ/5iicGyNUisYfEeiHm6tIen
wL3+p67DE0oHfV6S97a1q4h1sLZIBLBuzQzaLkbX8ZJtY1eXcRgOa5wjBqSkmjtR
sTq+nPIZiO+DSG+DzNVk3IkOJlwx6lM0NasXWSvbX1o9MpAPc2FUfqPYA+8N8s2S
DaO0PPuK2EKGDHtUSHzVd8tZ27yEeMJIRfl7u7sREGuXo/P0uPdSVp55OSuuOrj8
s3b+MCwmOct1Eib+9rxUKOs2xyGAx270uJ5ICn/VnOj1eJHAv8zpZ8+tTQXTZb1F
guFkM5GoUZkZgir3+950/Fc7AD0JQn5JYrIgCmaQMu9HvqaW0HaaTgYeC6jY2ViX
pf8ymjRu0Ibl2ePj0PJvugXpNYKtAE67NpgwiU7BijFBMN8XKttJt+1Ch4Rv7rYP
faP8pmOePBTkaakXDBb6VD8Zo6ta+19TyY2ZzoXdHJYhNP1enh4djaOWe1Yk7enx
7hIeOrAWbd6/j1/oEEW6DjkfrMMTM7Uo157qQDvvm7FlUdHY0lUADehwv1I3rrkN
1jd3lfI/QxJJPBeZKXxSWufgxvLi0bL///uXFe0oSKlQO4zr/bk7Ats3FWXw4+kF
0UdXnIVD+nRdLbTNx1WecHt28XC2pTlt1vyuMTcQF36/4s8+jRV52osVctMlQzGM
NdAzwoigwQ5y/V6yq4I3bq5Skqj0hVH/Mu8cOjVw5UHHtNgGWjcuzF0RaIa8TL8C
bV3PZZ0kRAPZ+XJPDc0Z4HFsFnxlgEFimG4Dikn3sFh3b45QuIwsoMvoCVUrjYjT
h3rfoXITv4xAo/5s4p+2ixGqOj8Xe819riDZElPrtKpeVutlHtRHxMe0hF48x7Jw
TB34/osK6MXlzX6zhVxxQ24IndNesNcvjoGQBSuVq3k6ib349tuTjn9IkuFR9uty
MlexG6Gf0tzjHNHELotBqViZL7VWnE/d1jHjyE5CbVdIPD/DfUsEqM5/0Xnz7w9R
uJvJtfb2FXFH5jDDAQW+TRpxp0ny1G1KrCdvxe/XlzJDPmkIme8ksVDnwHSu0dF6
zOT3krSvflwxiegBCCfbJHQWEJNAOus4ztPiWb0Le0GmpDYZM8CeFtvOAvO+JHTn
zIJbBfLvisqUMS1iCn3/VmBXKoGog71aS03hiHgxz9DFNjJmqZ2HHCGTdB/Ufo6R
Okw/2uPtOX3v8gAry72uCHWtBhXq2eq1tU9KUbpTxPnpjYujMP6x4TTrEA1jRd+P
0XKVYr1FCX6cQE/2GP5h1yJhP849xhzmi8wZqFmZUefbIzmE2SHSOsZsylp5bStY
dSMfc2L67au/QT2Ov+crJGdmKBQdX4U8CiQ54pocHtzEJfUNRRSbZpMAzfWP/LQY
h7m+QFfkW6cpj5hmp4j86RCM1cUy4gSVQqPh0z7Cjb4fgsgr/P0AD/blg7QbzFKx
WH4APC92VB53uF4yjrBCQ9M8JRynGTRUksn1MvUTbqbXXlxYUAd0cvdXJJfK6Fv5
2zeiNe5K2yry7dF32f3gT5oZ9eg6F5QFewnOt744ODWWRBWe5Bo7Rpgn52x8as9z
3L3GwyXec8gU93mpwHEuuZOK4ToYCGTeUWbwzWtMFrjnb38EQRFuP6TTqva4cgQ1
xEHp/67AJsk77UvBtnvUSA74kbMBB0ZuF5ogIslje89/wSeWGyNzrhHawt/f3sPF
XYpiD9kRmahLUICkj/JnCUfD+ql7Vl1B6TUIrJqc9S8m0lBBCK0IgtUjWgDTJ5HZ
Udr6Xz+9PPtE/JyqRKV5TcJneSQBztgQcGZmlSrdCkWFwit3n9FNNvLZuvZ1vBrM
z7K23aH8BVW+EQFsopNe9fKz8Ii9pc6Nx0gmKc8X5IttgPwlCY9ITu9HtAm4TYo2
zSoBGRLHpwu9LiUjTsvmAsRx52nEdHU9E4m5XzRSbU3LjxSF9CCW3CJS4eujZAoD
X9SBkLeTvjz5LzxLsoxDz25O8KTxgUfZbQ1I/R1fJSe5UCjDZypAAxTFTWhcy7tL
O0tevb7SbfvJH99IOh7SPmu4Or8jgzgjjg/vVGsSIcTL62kPbdW+71B4LXBGNA5y
wT3G2kdiug+2znc2DDcQUjU7FL19jqDgBLlddLijMWbhaBc5isYfdInFU6O5ao8Q
lDpQAQ1bDnOM0SV54J3mKKFNh5T+cMOro4Wf+VU3L3Rvnu0s8mtG3OJvwSYzut/b
Ol/Aokuvyr96c3GdztFfS/7CmVdTCyWbO1Hd/HSKIurMTUWRt7LYXFHT4lALg1SD
DIQDy4DVlMsdbTukdWv7itpvqpjMQFJ40x3ml4d1UVKOT/YAjOn0AZoRDka7xJjt
zYZkkwFjvMRVOqxSk6tcdejGNHYEit7I/3opbE6apbaH3XO2UxrH1q+3wCgICQHt
RzYcth0Wq14zBb4WqI0MXOo5Iv4zr+UgpG9bo+BCXWLOjVNoPnQbVVu2iBKEpYDF
N/wRPfRVP06Rm4xIAkZP769lBcAoUUx8BV/D0PN/iCH+ZwLFhTLpgjsvj1D7EjRd
pIAqJrCkHgCaY0I2UAY/gwkaEf0GSEJiiuxNmpFoHjou3MtNjHh62ejLgMYW0Pac
nKbax83PuGyJN0IktpmswIPeynfCSNd31VwLGHRdhYgCJA04ZpPE4WEmeb7wx4HX
SApPolW6bY06G304KN+laTg5DKtaHp0wDxAt7gLOVyvAVGAYX2TBGgnseWV2u5eU
DfMyAcKL82tptkVcCtmLZ04ZCbfHGYHAkm7Jv9xS+Ua+DBZux5/TcTuCH2X2hz0/
YLpI2P0vM08jcFiNXiyX721CJX7iyQiJV6RoS3nmheaJxrmA7Q8OAYvUxBPcf0tc
VC3P6sDuqN74VZ7jY5UyBe0IgH4ZXSDiPmImPyDHT9TnAEo9UuQVR3WwLsdGTTmR
uIlVn7XDKClziwJdA218MSqxRx7FHPDtHS3U2cRXZSpbKD7NFFrC5AVEp0r4cIM7
aR/dFkYDo3OqANUBs3s4LBLSoAvTnDEIeM1th1VBQaoSUA+vmcnjwWvLApYgpEv8
mvl6FAGdfHv0bx3ubN3hyOhAEi3QEGGHCndixPyLIWrKe8d5f9pliyHkbl8gOM1y
p0E8LrDLFMuBxsJ+H/cLwjhccFdZoPfJfyHfdJyUOMclFlxqDcME8Eg6j3OSHPSz
1C5mExvz4WLOmxtu6IooUJOIZd9SIV8QJkSOPvMb/jg8NOGTYE81eVjXlsvGy1XH
MX1gBJ4z+wt3Q901p4Vglg/KcqSypno3qkC7ckTYFKt5HYT5FK/fb92o5MOVW6mQ
2zBQ39NssuibZbMO/GNRX+oZ3DDdEG4l1Sk9/nFT5k8ot3VmIi5YJMtFyfBxO8UC
bw2TYae4GMTYnG6gy29dsx3gI0hrVG+kgBLEf+z5Cu9MoJifAMb1s0B05uMwv/gB
MYHhtHFX9P6fvgMO20Fzlez0kF1BVIBTmmHxlEu1LA2CWfeloVKpZxleohyUBkiY
yw2Jwl3SFHIQXidqb3M+1n8LoZwFQIMGXNLKiY6GqdHmzbxyRWYA18xZVgsLLkpl
cSA5QriqroUYA2SrJKJLrZY0kbnu0uzE5X0x/rl9Rd3VX8kQXJM6mIwlfu8QvWcc
TG2AQmyBjLAeFScqOgc1sjrnq100GgqIQmyPRyrEM5kXIpdddnXhZyQ07cXoaAwi
L9uE2ZpSEQKeC5dM9goHUGoZ+TvaSJi9oAe2Df1E3qvinD+PKsrrz4xmoU1hUKtz
Tcf836cZ0fWtNdZ4aENSpSlSduLOuAar52Gj1GaXYAAT3NC27fvrXW6hlWMAc7Ys
EYlgpnWG95a8r4bediQNKYjtGdTJxqchbdGCWZHtVo96Iha1rMxZsITaRe0u4UDQ
+D+ZQB1lNbjeOOQCGzK0Onbr5kPc5Wp37Fn3fOkcMojnwr8UY4CFMs33ZA42Ij4x
ij4dYvuAeNTeDvl3DeN9O3WJSq+FoudKD5j2RlaujsPP2iSgh42fqRnwvpNlfTRx
X4WrrG6lWe5x9W2wulHEz55QnlsB+d48DOAZQrxHtna2hB4/7DRjXJ403Zq9+hHX
MyZHzRaZGKpqUyHOvFQk00oie7JlmYQ1zFjkGlwvn5UAButOhcEJAYGBmpmyO/OV
2IvKj+bhMBLNr2HF1xnRaFZqJ+/E3T9P4pK+s2eSPQWGab173XP7rbeHZX90B7To
LqpTzzT8I/QVWA7k3rJTv2PGAduC7E3G0+qwuTsPoTvef9xpWbPe76eb2+rlVO8k
3ADLljMcVmy22JOrry/pEmfkh5dig27OarIpJxpSmcY4oGAipWraY8ZqfGZuHxPD
xdbbC5YH0ilrBgTdOn465WEBCXk5jZosfQ+XZatDMEtSH3ljuNoYE7PL4UcnixAN
GW9/maql25fRgpE97RYS3iaBDmF2dugpgwyurnoqY51wJOAuqSY1c5dTUNLR4rZt
vu3mEtnfpL1/gjRaFh1fzN90DjcKL9TdkoWCb2480xY05/7zdlrcNQwN+lx45Gz5
xtn+LnKiHagAOQO9BpHhVu9r5N2Ikbhkm/xXY0TdHU4ADwvWVbqvBdIijcx6/bAs
0yHUukvZYYmoxcahKtY+TgfVHaTfZNAGXiOGN8i3kewq7dB0qWv15A8V6fxhc/vx
8Mcm9U7NnL3LKsWi1fcSSKX68vpMCid4Qk0Od83BUFbr31ByLQD+6N+4dT8t79/Y
v864qHnGCxsBEK6/qN4DbBqYZpwB+kxRLG2qOGPiwUwkzQ3E7DL9cC3T1Pi74ypE
Xil7nVP6azKlSVAX10741y33AbCgLNUTlocS43lF7rIEBl2rKsW5nZkxzL8knx+Q
LHDRYJFrtMYNh51cj0URjebjjEHrwR0YSPQl4l+8Sr3rboBUym2WR1DYTm4YBKG6
8/fJwyZtBxZS9/fW/lC3IzLX+d4KC+Y5n+ASrqk10ZsQjW+zlVi58nclsU1yBs8F
PKvYpetqT969tpeSIpe6GBVxQzCMQPD9N8yNMcpUXHTwa77Qkh3LHQY4KAWuyiMw
GEyZZiBF0wRO26aEWLZLR6eF9gFCcwxEMhYp1X2i8Z4NPf7QAgNDBAtromcEF3sQ
ZEzJiHBFGiBrUxNMC9fcqFA9sJs7aYBzbtuVq56McKWfzpG5IQlzWD8TVKKeXBOf
iM6sfxMD/85iOHvLMj27HPlNdJc9MLqOjSJh/OK3kmQnuP80mdVsXuGTsNeA+HY2
NPOmhIBK72MSlX8Xj8sCc5nkG9AQFh62rgQ3MKu+KrRi3MJQIVqhuOCwOVY3Nynx
D8fGpMsEWkvNmmgP0pviJDg55LtUc2xBtWMb4z18MGfuveiQdiAUo6WyLC2nCBg5
znzv/BBkDly0TECCYZ/5mHVhduoIdxpzQZrogWCE8JcIPofK+vwx/ztRAdla72tw
/GZty0BX/xelDl9nX3imRdWlaQlaQ30s3Z5+U05Im2eJLYK3Hf8ZDYeDn30pMEIw
iREP5+lrA8wa342MJQQ379SvIfRLHFrqol/4Tae91TjEJUfJ5F5L4SEG9jKCGNwe
quhxQk8VvEpDl0ggkcfaXB+2IALcIo/ehSIpqXcAUgsnaGJRl+xHxLme+Ed96jIa
X+IvhKnoAcadIBLmknJR3gOvO+AeFSU9Yq96QAKKAVn5Wgdb+5HWHCQjfyxbBaBv
5z5MazaVigjfS54a53aLpPC6usVPGCXKeffTqPh97XIR7DEmSSW40FpGXUnxXFPX
PVWyOcdCBy6OpRTYJTDBbXGDaTk1sphNHe5RkR948Mo2k54GmhibCwWca2r1SBNW
QOyzK3NIJPFzx6VQCB/0Lv1yHMd7NEXdu6XlFhAXW3FvXYH8y2sV25Z0FI3RWsOw
84Mz3aThDJIpnZ27SWA7uoRnjWrMznydTseNBhgJApce/7Go8IcYUq7kOCJ16+Y1
L86Jo1A5rECgMyH7qhuE64fkKk7tV+iBT5JuSb7nrnvXL7VGq7qgZ4eMH/+FcyvR
edQpK+Pi+XxF/YB9RNQYSf38dYBue3U3f3J0bpfl02/pZJkrlE/fmoP9FRHaog9v
t8wGXifA4bJN66Y0/b+jSLFC6qJyJDrypgNWN/nHbI7hCyUSHc/PauGsTYlcu1B8
CPwZdwtcCpbqadxbiv9Kaiuyxv+njM4qhErS0wIoyBYm5xbIYV67KElz16Kxpkw4
EsDV74PrJE1Uz5lPm7gAtPIyNh+mRv2FWbiA2Jj3dVe4bIAvWmZ10Tavm1Ysyb+Q
s2vY6QlFnlC2fF/MDndGEwfDliAUfKaIG1YzffdBEtYhmsSnR8ZMve5JnohAly4q
4cBJI66MEP+nc1vJqAgk88C3stUnmUJSCmAetbz+FjPB84q1mq2FqfmoAAG93S6g
slXzhTPtVPm8a1D7lGvIRVNSkpnCGMk2iC5lUh8g5xwPuqoPtX3GIiYbCdAJ9eyt
JNSpNQcEyIIU5hvr7aX7X02P55BAzXet+0XRZ/wxg0+KpyzTwkzc7fv1YDO4wW48
bOYKqB/CDJ9loJ9fUuVPKqefwOVtdpUWmslT6SxVZaQj9qQJwrC1+p5TDyK9zkhI
9Y78PQwxjpwJFuEH80a8PPfaPaosOK24bSCYsvExLpWnbACCLKPGg8dgEEY9aDav
oTtv1tjhtcogQCDUaQ2jz90+so26NopW8pfyC97JVFtYBORF7K7W2uaUb+Gf9KuH
Ve1IdqfRGUbEQGCASYQvsCdW52ShUdBqPXIjxSps1kPfei10JzUj2mmhBfy3HGAj
S6YipHLEwRs4OsX7nvHestS4G7gMyOlsu5AKWHsrvW6wO78As0noiXG26EO6Mdic
u/LAVk+ie7vp1asr/RF8EEvcRRSWIdCkR9QEuHrvLNtGSct3qzoOj6gX1VcuAII+
+Do5RGk42qJKbhjlFvyaK4ccKt3EJ2Vjj2lumlTxzfnDH8Z7yZJrOvgc0sEFEcwF
kn/xaK/hC72BS1zJcRqqmP0CiXA859REt2u9HDwxSBTht2zhxwW3VW4WegC+9+1g
//2SnZJCsVm+2E/tI/pjnFjQvGw6lZbsvwOXhkgMcxGbcx0qIahoaIrXzGKvOiHz
rnqJEUbGb2G9VHLNNRcdEROu/9OvuYLESENrEZI0n8sHqPig/qwbQovzzViMZ/DL
IxShDHnXDQMNVGpaklK5fpLX4WIO2r81ykqh56y5P0xGMHPg5uAgw0lRfA0qz2zQ
Mv1R4ZJuxAg3MjDhs3ngKZaWNFSEauIYyQlN+6mpO6UqCtzdDC8gVs7kMU0BH+o6
ljnMym/FhjYb752L/rYEDztbHRLzFCd/eGgJ52acfETrbJaVXSPOho6KjD+R9lnS
0GiBxLqvSwmb83js/wo9zQNu12Vi4W/cAs58uKcK1UP6rGzct3SMB/60kjHzsfU1
g0W8v5lX8/DkUO4oWXHJmIoAliCUqRhwu10WRrQQiDSJPKXS+qerBVJTokJJLE74
NWNSIX//lDNNHVWGs9AXgA==
`pragma protect end_protected
