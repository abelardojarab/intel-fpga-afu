// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// Generate one pulse every 'd81920='h14000 cycles.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_metronome81920_3inCtl 
  #(
    parameter SIM_EMULATE = 1'b0,
    parameter FEC_AM_BITS = 6
   ) 
   (
	clk, 
	sit0, 
	sit1, 
	plas, 
        sclr,
	real_sump1,
	dout,
	reach32
);

	input clk; 
	input sit0; 
	input sit1; 
	input plas; 
        input sclr;
	output [16:0] real_sump1;
	output dout;
	output reach32;


reg [16:0] sclrin = 17'b0;
reg [16:0] ripin = 17'b0;
reg [16:0] sum = 17'b0;

wire [16:0] sum_w;
wire [15:0] car_w;

reg sclr_r = 1'b0;


wire  [16:0] sum_w_1 = plas ? sum_w :
                       sit0 ? 17'h1fffe :
                       sit1 ? 17'h1fffd : sum_w;
                     //sit0 ? 17'd32766 :
                     //sit1 ? 17'd32765 : sum_w;


wire  [16:0] car_w_1 = plas ? car_w :
                       sit0 ? 17'd1 :
                       sit1 ? 17'd2 : car_w;
                     //sit0 ? 17'd1 :
                     //sit1 ? 17'd2 : car_w;


always @(posedge clk) begin
//    ripin <= {car_w[13:0],1'b1};
//    ripin <= {car_w_1[13:0],1'b1};
    ripin <= {car_w_1[15:0],1'b1};
end

always @(posedge clk) begin
//    sclrin <= {sclrin[13:0],sclr_r};
    sclrin <= {sclrin[15:0],sclr_r};
end

always @(posedge clk) begin
  if (sclr_r)	sum <= 17'b0;
  else		sum <= sum_w_1;
//    sum <= sum_w;
end

alt_e100s10_lut6 s0 (
    .din({sum[0],ripin[0],sclrin[0],3'h0}),
    .dout(sum_w[0])
);
defparam s0 .MASK = 64'h000000ff00ff0000;
defparam s0 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c0 (
    .din({sum[0],ripin[0],4'h0}),
    .dout(car_w[0])
);
defparam c0 .MASK = 64'hffff000000000000;
defparam c0 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s1 (
    .din({sum[1],ripin[1],sclrin[1],3'h0}),
    .dout(sum_w[1])
);
defparam s1 .MASK = 64'h000000ff00ff0000;
defparam s1 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c1 (
    .din({sum[1],ripin[1],4'h0}),
    .dout(car_w[1])
);
defparam c1 .MASK = 64'hffff000000000000;
defparam c1 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s2 (
    .din({sum[2],ripin[2],sclrin[2],3'h0}),
    .dout(sum_w[2])
);
defparam s2 .MASK = 64'h000000ff00ff0000;
defparam s2 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c2 (
    .din({sum[2],ripin[2],4'h0}),
    .dout(car_w[2])
);
defparam c2 .MASK = 64'hffff000000000000;
defparam c2 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s3 (
    .din({sum[3],ripin[3],sclrin[3],3'h0}),
    .dout(sum_w[3])
);
defparam s3 .MASK = 64'h000000ff00ff0000;
defparam s3 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c3 (
    .din({sum[3],ripin[3],4'h0}),
    .dout(car_w[3])
);
defparam c3 .MASK = 64'hffff000000000000;
defparam c3 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s4 (
    .din({sum[4],ripin[4],sclrin[4],3'h0}),
    .dout(sum_w[4])
);
defparam s4 .MASK = 64'h000000ff00ff0000;
defparam s4 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c4 (
    .din({sum[4],ripin[4],4'h0}),
    .dout(car_w[4])
);
defparam c4 .MASK = 64'hffff000000000000;
defparam c4 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s5 (
    .din({sum[5],ripin[5],sclrin[5],3'h0}),
    .dout(sum_w[5])
);
defparam s5 .MASK = 64'h000000ff00ff0000;
defparam s5 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c5 (
    .din({sum[5],ripin[5],4'h0}),
    .dout(car_w[5])
);
defparam c5 .MASK = 64'hffff000000000000;
defparam c5 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s6 (
    .din({sum[6],ripin[6],sclrin[6],3'h0}),
    .dout(sum_w[6])
);
defparam s6 .MASK = 64'h000000ff00ff0000;
defparam s6 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c6 (
    .din({sum[6],ripin[6],4'h0}),
    .dout(car_w[6])
);
defparam c6 .MASK = 64'hffff000000000000;
defparam c6 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s7 (
    .din({sum[7],ripin[7],sclrin[7],3'h0}),
    .dout(sum_w[7])
);
defparam s7 .MASK = 64'h000000ff00ff0000;
defparam s7 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c7 (
    .din({sum[7],ripin[7],4'h0}),
    .dout(car_w[7])
);
defparam c7 .MASK = 64'hffff000000000000;
defparam c7 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s8 (
    .din({sum[8],ripin[8],sclrin[8],3'h0}),
    .dout(sum_w[8])
);
defparam s8 .MASK = 64'h000000ff00ff0000;
defparam s8 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c8 (
    .din({sum[8],ripin[8],4'h0}),
    .dout(car_w[8])
);
defparam c8 .MASK = 64'hffff000000000000;
defparam c8 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s9 (
    .din({sum[9],ripin[9],sclrin[9],3'h0}),
    .dout(sum_w[9])
);
defparam s9 .MASK = 64'h000000ff00ff0000;
defparam s9 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c9 (
    .din({sum[9],ripin[9],4'h0}),
    .dout(car_w[9])
);
defparam c9 .MASK = 64'hffff000000000000;
defparam c9 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s10 (
    .din({sum[10],ripin[10],sclrin[10],3'h0}),
    .dout(sum_w[10])
);
defparam s10 .MASK = 64'h000000ff00ff0000;
defparam s10 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c10 (
    .din({sum[10],ripin[10],4'h0}),
    .dout(car_w[10])
);
defparam c10 .MASK = 64'hffff000000000000;
defparam c10 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s11 (
    .din({sum[11],ripin[11],sclrin[11],3'h0}),
    .dout(sum_w[11])
);
defparam s11 .MASK = 64'h000000ff00ff0000;
defparam s11 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c11 (
    .din({sum[11],ripin[11],4'h0}),
    .dout(car_w[11])
);
defparam c11 .MASK = 64'hffff000000000000;
defparam c11 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s12 (
    .din({sum[12],ripin[12],sclrin[12],3'h0}),
    .dout(sum_w[12])
);
defparam s12 .MASK = 64'h000000ff00ff0000;
defparam s12 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c12 (
    .din({sum[12],ripin[12],4'h0}),
    .dout(car_w[12])
);
defparam c12 .MASK = 64'hffff000000000000;
defparam c12 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s13 (
    .din({sum[13],ripin[13],sclrin[13],3'h0}),
    .dout(sum_w[13])
);
defparam s13 .MASK = 64'h000000ff00ff0000;
defparam s13 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c13 (
    .din({sum[13],ripin[13],4'h0}),
    .dout(car_w[13])
);
defparam c13 .MASK = 64'hffff000000000000;
defparam c13 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 s14 (
    .din({sum[14],ripin[14],sclrin[14],3'h0}),
    .dout(sum_w[14])
);
defparam s14 .MASK = 64'h000000ff00ff0000;
defparam s14 .SIM_EMULATE = SIM_EMULATE;
//===================
alt_e100s10_lut6 c14 (
    .din({sum[14],ripin[14],4'h0}),
    .dout(car_w[14])
);
defparam c14 .MASK = 64'hffff000000000000;
defparam c14 .SIM_EMULATE = SIM_EMULATE;
//----
alt_e100s10_lut6 s15 (
    .din({sum[15],ripin[15],sclrin[15],3'h0}),
    .dout(sum_w[15])
);
defparam s15 .MASK = 64'h000000ff00ff0000;
defparam s15 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_lut6 c15 (
    .din({sum[15],ripin[15],4'h0}),
    .dout(car_w[15])
);
defparam c15 .MASK = 64'hffff000000000000;
defparam c15 .SIM_EMULATE = SIM_EMULATE;

//----
alt_e100s10_lut6 s16 (
    .din({sum[16],ripin[16],sclrin[16],3'h0}),
    .dout(sum_w[16])
);
defparam s16 .MASK = 64'h000000ff00ff0000;
defparam s16 .SIM_EMULATE = SIM_EMULATE;


wire eq_sclr;
alt_e100s10_eqc17h13ffbt2 cmp0 (
    .clk(clk),
    .din(sum),
    .dout(eq_sclr)
);
defparam cmp0 .SIM_EMULATE = SIM_EMULATE;
//wire   eq_sclr_short = (real_sump1==17'h147); //A10:'h149-2='h147,S10:'h13f-2='h13d
wire   eq_sclr_short =  (real_sump1==17'h13d); //A10:'h149-2='h147,S10:'h13f-2='h13d
//wire   eq_sclr_short =  (real_sump1==17'd2560); //A10:'h149-2='h147,S10:'h13f-2='h13d, Faisal:2560
wire   eq_sclr_0     =  (FEC_AM_BITS==6) ? eq_sclr_short : eq_sclr;

wire eq_sclr127;
alt_e100s10_eqc17h0007ft2 cmp1 (
    .clk(clk),
    .din(sum),
    .dout(eq_sclr127)
);
defparam cmp1 .SIM_EMULATE = SIM_EMULATE;

always @(posedge clk) sclr_r <= eq_sclr_0 | sclr;
assign dout = sclr_r;

reg        sclr_r32;
always @(posedge clk) sclr_r32 <= eq_sclr127;
assign reach32 = sclr_r32;


//==========================================================
//==========================================================
//==========================================================
wire [16:0] real_sum =  {car_w_1[15:0],1'b0} + sum_w_1[16:0];
reg  [16:0] real_sump1;
reg  [16:0] cnt1;
always @(posedge clk) real_sump1 <= real_sum;
//==========================================================
/*
reg sclrb;
always @(posedge clk ) begin
     sclrb <= sclr;
     end

always @(posedge clk ) begin
     if (sclrb == 1)
     cnt1 <= 0;
     else
     cnt1 <= cnt1 + 1;
     end

wire   wrong_0 = cnt1[16:0]!=real_sum[16:0];
*/
endmodule

