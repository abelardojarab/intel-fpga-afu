// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// 8:1 MUX of 1 bit words.  Latency 2.  Select latency 1.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_mux8w1t2s1 #(
    parameter SIM_EMULATE = 1'b0
) (
    input clk,
    input [7:0] din,
    input [2:0] sel,
    output dout
);

wire [1:0] head_din;
wire head_sel = sel[2];

alt_e100s10_mux4w1t1s1 mx0 (
    .clk(clk),
    .din(din[3:0]),
    .sel(sel[1:0]),
    .dout(head_din[0:0])
);
defparam mx0 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_mux4w1t1s1 mx1 (
    .clk(clk),
    .din(din[7:4]),
    .sel(sel[1:0]),
    .dout(head_din[1:1])
);
defparam mx1 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_mux2w1t1s2 mx2 (
    .clk(clk),
    .din(head_din),
    .sel(head_sel),
    .dout(dout)
);
defparam mx2 .SIM_EMULATE = SIM_EMULATE;

endmodule

