`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
G19eJEdTFa7Sn2UKlO1E0kN9e7qzsV3TVxSQM9QBYgboURTxrX3KvAQpXFk3TMD3
/CS9lBQ0jcC5DWut41AwAaCMdIBpYneC3zRMbzByOLvlXqop5E0hBNrjThm1K8Yg
5ZZ3GR9GjTdmgyD/lIMSlobxqXwNVer+3Qb1FLWmMv0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2992)
tofqNeSfNIBr7+ah3l1cYOS3spZTcYKQfCUgOKdhLbTjldWOqDVHao7/LhpxgbLG
zbsiu0FfDdtP+BDA4sQYlk6iysZuz6XtIPMb7pW6P7+7sksq4JDH6VA83OipBZwr
TdkNOHcJUTTFkECRMhsVW6Gv3MnLvY5ZP7RkZa2Lf/G8NDYkP2SBGJZUd3kMRVW5
wjdYEMK2HRJNSJyOX046TUhPCmIge4tc50ZojP92u/0f+qlhoKSU+dsI2c5UWf96
F6c8w6UGtrJNTZCFJBxIVYvzV32gZwi9feNz4Q1ElHFHtXtjG/tAUp9AOpXTndSD
vN09oVWHVfavqodepbD1v6Iur+fdyNto4gMoPOmMHcp8mErQv+h2AqmvFdPkdgxd
ZgWfI5mvOUkmgqV48fVV0ojo95SFycZg1LxUuVh+sjMhhdcLMWmUH6/ycg4yvOKZ
iott5gx08xm4SauJuX8aV5+hno6DIRkPZ6xxM6F3I1JWR9+r5doypftYOuaVelIm
EfUeMmcJKoPrV+u/kYT1873Xgap9UuIJgvYL3ritVRh4gcCx1q3TFKuktKBIhiLA
TZF8vL76LDOt6KG2i1NBRRy4R9TZReu168/0Zg/6oiJN+FGGXOgT+g1HvcCgKtlg
PLgefb5cNmBVE3EfR/M1UuxFFPZIIYRSFe214I7JIwH6yeW39n/VIMK5hVzQxPWm
KVmqMofJZtDNqTrDHgY56fN36nUq3nJC7tpGxDlgDlth39O92xvqxEDvCKNhhs94
FSpblCASjzUM2no4SFPQ2+E9ZIvMbzhvDinbhVt0gFOZQRBrJxS/6nc6GLrUjtt1
s6e3WZ09ch/iiBAKNh1mfwixjfONS2efpRCm9vdNVAzocinqD8V6CnbngsOqJIkX
0fQiLBARDnC7BJ9CF+qiYLI1WBbR133jrYAnvkaTJOJyj28JmA9m4yempCJ/pG/D
KzsCbReXtmt9B6BqRBBnj2QeCZ99npzzlQZET8VfJy1oDLzT97m8iofL1oXdPcuu
1WtsLjlFuT+TzcmYUkLmk59CbWpCgbM8TwxZajdyubg68FfodF2SaiEFyQ+keM72
FNK6BzI+ELSa3dzeqKOWS5oW+ssJ0CxQA8JFtadL4LFyYYshvVGYebbf+N4mXdII
coGz0KKoJTZpKU5WxjrNXrY0OEBeG1/ufzaZeB8Idr6XEqRAQkbgCXX03zyOEudN
Z3jq2V+NyYVpcdejCKZzN4bsp4IEWQ27xsCHS9UfAW+g4stsvnDrOX67ZMir+Jez
agyBFUUAdJn5S9vNGSfe+KErhdT1W/7+eQVSAbizO6H5HAjeK9Y1xUe4h587nUQp
0C2zjq2id3KkTenuj84ilOB34g4BnIonff4KywKII77j87k6LwkzbJPSBjbnHfR/
FA9jfLMhgc/PHkfDKvxjbVRTpHUlLfXMm/v4QFUFySgDy5ei+RbpEYKQc350fGJt
di8vhQ7L5BI36pVWsNMRnIy5H2Yc0Ftusf72DtPFiUbZ19D1GXCKuM9B9lLDhltG
14CQtjxaFG17h34mjNNV2spihq9zvv2OoqopQcPhd5BpK7yVKPbAXU39PN3rQaN9
DxqO9Ze7v+g/m52/c0KAgQfiZ4Buv5cFTeU3e6Pb2uTfB7hfgKAjyB4yAZkMTLyo
B6hZ+am6/X0WsrB2zPtce5cjDiFhcBbNGvpbbIFmQcfBTeVEiFnYUVqQhwYwjaiy
e9pQl8vVdE/q+FEErpOouC9aQd4S6p50blhnsQe4mQBd6i908SQ4gbxzwQ/PCRCT
nvR/S4mzjbr0TWhjtZDZr6XtlVSLP2U6DwWDRZz3Mz3R+3ftUeboEK1uM1s3p0zP
CORZGjg5ZtIgxXmi8tWpC7AmPc+Li0JdGiJTHPmtxftpogub/dGLAbc4twDxm1g9
shgk/l5S5OLH2RGnK/WQBzqOLtclWiLHa47DnRP/zR92/vH1kJLR2Cz7YmRVduqs
CvW7AAUAodkswG1P2XAcsv5SGAEQUybz8it4umCUis9K9pCWv37DpJCmE0J9HpLx
IMc7qdid3nTHXnw7dY/Gyq/Useyaay4ItPQoCDN6VZ+fW/QuMe6EwcYhluCN1S2y
237mGs1iCB/HGmI8l5eKPjm8DTeZiVA8Zb/pC5OF7gZ/IyeKCTteZLXrEbScFcLT
x6j9yLGH13V2sXYK62vuDOZYvYatvpQLsi6Dy7NvDmu+XGobEjrlF4cXxk4swRk+
4j2Aw8MywthYelqkE4X2rkjaQ7Oqq5m2mTKl9e0Wy8+/klv4WL+zPi32VdIjmtux
z5QkH+REk+UGs0ixNmlWTjbgE/FQyyMVWyjtz0uHbfOouxB2N8yrY/AomGJp+VTW
S4JVsQOmtO+dNPF/r64pqURKazY9Xh8qyiGFoeyJVAVb34zC/BWq+pnaTICqGv0+
ieKhSL4cvfvPtGg0YPOH9nUdGDsfrLj8vSD5fkZBgoPhiEXYiCmqsJqjloh7m2h+
pH8YOT6r9ooYwKGC42jE15+7bzZV5wAmV8Fb3bjREYMcIHPkEbrqJavGICjAjHWi
o5ya0t51nLMuludS3hfsX2hvqpQzkqa795yugaV7cNRUpNwGc7WaLfsC71hK+5pf
uy6zlCDJXu+6/tjPiykDfLoK579EjfYdKmYUSeYz/YoQq2k5d9goXYhKstpjfA7I
98LcgsSQpJXiKj26rhOb5auJ2kRT/+L6LJ1d/E0JZ1xWGFK/FF/mwfl4wxL2KMob
HkU477p7twajtXTux/FBcT8UEEd//IqDDtQlehU9uK6LYFSESk+/vsYC0pWnSrxd
yaKvQ3tiNgirQhBUWmSAqRdonu0JKu9EPXTa9BVYCK9H7K3c06KwLRmLkLKhhivn
mtNaJiY82TA0RaVUSD38ZKsAbAk0BCvtpBcJWv//EDaaX9gs/yhjW/rsqEeB18Qe
f7VL1MXZgoCXJrCMmQjbu3EW9AJfQZaCVWzHT+4jiPDlCuLDHReKin6yckS+QFzz
1l7UT1shtY4GpCARZh9onaDpg8PYa/r8B3UVufGb2FBATKykl5n5MPxRLEfIW1Pd
P+aF+YNnCY4VFz+4SMQWsfblq98gsjh1hONzOAq4ObdxdzIsWHOljKdUIlW10e9Q
F3Ue2m9ZHNu4cJvozkrH2yzDhyc1BtBhqWTFKpeE3bqgOgG3quTIQwS1rfcE51xX
dEQgZUqmLMThTKZZfxv8gj6dZXmQgDvetT0XdLfOS2vcryYkYZjNGyj7vdHp21ER
TdNEewXTG/sETAc9UWyj0FI7Z01D/ZVDkbWx/Ty9YABjLPNBIeaIJa4Sq6oYQqrt
tfgu9L0TFX9n2/12WxacDidiaU6QIUrPNmQWdqtUY+0yPmlRG4gJV5gUXBp/RPL1
ddtJLvt7G9Xn+qb2KEdPlfo670ELyfqC1PRL5xnrXxiYNho5srwr+NUvtHVIg1zJ
durHo0xmWmmm4sUd8qEMWUlOjo0qxSs0TiV47qef8FLXuU/bvF33mRlPUpHyyzR+
V40ykajVQ2BrkfQW1wikPbOxltPPlnuQUSOueIWgopi1WTAt4UBwkh1Kqhi9z9Jm
PYgaqQ+32YsMtyQGSKzNTne8yK/9M6SELIQl+GUzaaA7nRzacLg04n0Pm45IV70t
YjY6jQQ1oWUpzM0ZrS2x/WIzRzPGV949LEEHh5hzEVG/x87PCJgzeGpJmV4WKjXy
EUpL/Nt+JBJHqdrZBCnFOxEXOCPiXg7iEcNoiZrR2zuIn/YoagDHqqBegoQ/HJr3
urfWitAZvbke1ZdJsje3eHYSue1R1Tdm40N8IdvSyulaRFvzDVpFHrX4MXWLpFUo
vzjkTDWv8wJUbBsBvRiryCU2iLB3EGfl8O8z/3iCLjj1WairFfi4shxG/EWZo5AW
U/ASnC7wmO3xjJ4bfinloNI4KIebWsEnVY0BHMPuqm7svYuDNj71rGFkLmKTaFMh
Eqch+1bwmEIdc+kqcyKheA==
`pragma protect end_protected
