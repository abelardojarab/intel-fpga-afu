// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// 17 bit val == const(13fff) equality comparator.  Latency 2.
// Generated by one of Gregg's toys.   Share And Enjoy.

// 17'h13ffe = 'd81918
// 17'h13fff = 'd81919
module alt_e100s10_eqc17h13ffbt2 #( 
    parameter SIM_EMULATE = 1'b0
) (
    input clk,
    input [16:0] din,
    output dout
);

wire [2:0] leaf;

alt_e100s10_eqc6h3bt1 cmp0 (
    .clk(clk),
    .din(din[5:0]),
    .dout(leaf[0])
);
defparam cmp0 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_eqc6h3ft1 cmp1 (
    .clk(clk),
    .din(din[11:6]),
    .dout(leaf[1])
);
defparam cmp1 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_eqc5h13t1 cmp2 (
    .clk(clk),
    .din(din[16:12]),
    .dout(leaf[2])
);
defparam cmp2 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_and3t1 c3 (
    .clk(clk),
    .din(leaf),
    .dout(dout)
);
defparam c3 .SIM_EMULATE = SIM_EMULATE;

endmodule

