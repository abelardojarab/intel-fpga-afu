`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WtN6dOz7H7bxL92hP9DWuWj1A1tTv4xq2TZBbEOT/Wca52eAGvrpNP/pTC3BY8DV
RCF4X93q3quYagQ5dQjdCDq/5ia1IjHg+WeoZkG1cMzXGYHpgiNlYwbkVp3/Ku4d
GLV/64X2ZO4r/YvzmGXhbbip6lGZeiQO3I75MXqe/+U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5664)
u0BDc3ji6LBZufk+ioilgjA/bZSLlUazYvADddtCxKaSX4/6OHT9xXAdO4rG/WDF
DnTPfUjsmPw7996/wNxXKBm0T7Tn36qmrvjHHhTN+4yo63A2aMcO/EYNJaAepAAC
m+5/C8jBP51BRo2UmBPDzXBXOlEq+yfYnlqY+l9J/EFJZMvF8Am0svHxo/k/bjGE
fE09Zs7ijbFbFFYA7Z7RAuVWkWSWa28leE0yx1Ffu8iLufPplNrl5oEkDLJCad1A
hwkQhTRM5CIG8aMkCgCn8KuV9ezl31JcpyLpV77iUFlNlAO5QolWMjTDcf55CIWY
v2p6BOwX1wSYloKG4r0oRKhmXmJbJepfRS7M7DCMdQ9cLk74OunqIEBBDwACpU9S
Q/BSaZo4YESrfRwNcWLNJOqxmMiKu1zG9qoYOLFV4+wOx/tNzSYTS7UpBL5gmaLP
su8RuEpafT9CUMacbvU94/CiN9A3Hv2XGtpN1ovIyFf5SiQxVhWjfSxSqJsgTnVK
iJeibq/+VApfUhQvUE0WRkwsA/rCml4FXI1zUKNOckmUMLcKCNuxzKSbAW4mM78y
FJ5FY5VspoVd1lTVvW14B1WGKiseM7+R4enBLz1ROSInHMHzBRR0oex+gR3hpAy+
hWRDOCXbdmXrwJhPdFTZeNw5xunNAA594U7Hzrzp4Xt9l9UxAQNwmFWDGcGWga+L
u1z9HlgjvEjVnl513XrsITu2gry6nJsUbBAuTtUkJqktjIVp3L7qvmUSbM7QlNcu
v4nmCajTx0uxRLC3JLZ26XNOqj99KE2drkUb3705oLHQ1Zqb+I9LzJfOvacA12hd
AOQfhR9dULPk3RWlCyATrlyxuImNgv/nzZJdr1sm49ikxLZE0wF/pT36xne4ShIJ
o+YaOF9llgHeruSFEy3dRD4rNziwsuc8CBGCvw430JIYKyXSflci4W/YnVLYinov
h/JkJYeCi9DNwNH7Yu9gQvXxsCcp7kYPmmGjuIk6qLmg4zRwZCJgES9TsV2LSsDT
nYeJ23UlgrA/fJbZ+fAAv2WtiJh6K1jvqeYDDkDRKSiqobs+o6/w7TqCcy3xHy2m
ZWaO695XR1GcXRVSWrNOhV+uEUhLSHJRWvqX6cndrN3pooyQcSU/CwISS8KmLFqV
f6nlRai4Dg2Cem2/Bdcc9yQZBkN2eGHt9189/CgCc7SOB8mtkB95dsQd2C/vCN9I
XTqoSAG4pq9XnBQPslHhkfoX5kDUEOPtudoT2250SrJ8YWnVnYDQGtw5ugnpt3ei
u4qr87tJnJ4rMrJVnzmHv7uDe0oru7g9462OCldUbOgHg3PPGMZv4hjhaciNF03K
zznrwI4RsDfa77KOXAcxqwUpkFqizh23vW+vBMFk7s1D0crywt3f0Vn2epUtIyda
mHIoAN0WDB7lX5jhaBg4HirTS2MXGo2SHOaIFsogiz0XHev0rgcKPC5ZrjEkRaeY
NJKuyvZZexLnkaV5hhVwjcBv39B8GP++dHftuiVlw83eVgeImpUoyWp6d8ljNxFN
QH4eKvYeL4kQGK2yld6OTNFeztcqKyk5eJfNGzKDzwI0Hkp7UqoANhcGurYGtQs+
/ZGLWD/hL1UvJwvXw6tUwiL9XWVfBnnI6UzyFA6wwWJ5hPtQO+ega9+XgAfZU04S
qyOZGQUgicODUlcPbQ1yPDJ9yLIPLorEe/bTU2Oy5/bTTcDdTkp/JFnRaVkgt74y
kXZ6nqKUNOB1VI1vsm2xeOqvyWx2xk2cEYsbt5SDMEDlP7R1ZSUtIbjQxwWqnYcP
B1aEMUgFHfOpbalVvnfLJkbCUwrksJ0IH1qtyooG2zPYbhdxFyIkcHq5pw4fzqu1
IeD900nxgI6KXrvoEglGNnYW3phZOzhm063JTOi6pPx20VE8h2g5HtiAIr6/OiNg
1fmPsokPfU/eO2X6frhGf2bBqaFVLqQiNZAiD6gVrzmVOLQMFJHDhQ+ZgR7XoD1C
f6uxSjx+IGkDt306F+ztE3i+WvWoALUtZFS5jAe6YeSW21QG+1nvsoXazEIIFJq/
bEidXBsCex7LTsnTbLY4CRbggUo6xHtXFCSp9XqRlcpnDq29KEQikXKJeMQV0OiS
zP5KyWiii1X4iOM2CBpIsS7HOg5Vf1tH2W6th85acufTk0eYcv6INWqsdJaDGwBB
crJ4XKM423ib78ExqIWVDhsE4am54pjBz6HZfiVupKxTwnKrVfNiYx99X4SkNR1m
e5+SQFyToICeESWfwCYqpeEAAvQ88PiAjl4CAf3FHEs7WlhwZSu2Wvfr/J4ugpjI
9tZM+Wym49bkOnRwyT0DBDgK3S7gHUDZddRgTKToh04LWQzdPxRACZ9McQDDNxQH
KUcwdpQi9NqH0npDFL7IqsU279+d0ufEGp12TqiSYkxgKR0Rm2K27K5a0D7jxv4/
of8qdD+Y3hnujEDIFtan59ERn8s6/8rKcmZ2Y3DF62Nsf+sFit0sSFej43aAR7n9
/baqfWFxO0G2Bp4WmYKkCe8vcKbYU/IM/UWwNwv2r1GlWMK87B76LWO96FRCOGLQ
TT2lQwWb7REYYrB8sJwGLjbM5fH34CEtpQk/IlW8S1XhVRY05HGwKT3Y37pkxPMx
VYc9WLy5IOsrgKjg/gERoOtyyvLFeyb2bE5j/rwbPIIYcwggYKdgWrp6kggVECTF
GOxxwjsYGd1MoZvIQP1mDUg+haX2HJL5xjDSCqji9DMq+bmMph6Ds1sdl6o3NcLk
9EB0IOl0Jhhpm1Xcw/Ecz2xY1JIOZPiqjsiVvmRndhZ/YWyWiPm6NEpDYardUYC1
G7vYnyKOWGcCL1xXgIKh06VgkgVgUBC/hw4yajwhWMnClZw052CL6NQPPudAvDlk
Hi5z3tZoilZql9KshSrKEYLHg7xnnMJZrmuC+YlK/xpWNy2hbZRnWVFtXm4r780w
i9Che879O9f4g806k7j5OeIczdQ302NXtOU0J2hC5r0ujDRDH5WGOiBHAYN867h+
+UslbUJMMYJv59pCD73Y4EEDNyG1yTSsxLFH3xKhTKCsuVilonOdLD3siQjmL0Me
HVzC1/gqNPnYMdoNJIuJ/cficVKDBBttZGi9atYjtcG1GWEKv81lXrWC78w48soa
NOwk3VttNtrSssUHtaJRDzbL1McK/NYU+8m2TpPjZV71mOOHu1yU625jjd5SVu1V
Egz7MdfcH/kixcq6HXwE3YmRhLzLw/BC2X5iwyS5TRmsNSMiGShiU5gIOgHCtVE1
FgKUwYIvrcq768ZiLldY8vwPOOFehqfVGsGZ3VTKzydyYecMwBCcgyIB5ZxxJRJo
sc1l0wgeH45081ZTjoEsdcUfdqbZaTxN7iJrYGFu/ItQ6QPDvMqQp97RQPmw7KdV
T/Kp574dmIOd8qqud8p2JEkN63UaAjCwYrcpraT6G8qT2WeKb1iuTQEQ+SWVj411
cGF+/oPhumZKOvfyA+4oCRyI8OmPHAywXuMQG+HA5s66G4MaXGvyLdZC2QiVDzuQ
l7I1A/sAJX3D/2d7GlQMgwiOYA+lWZq66KpOUJt+6mZyGItG5zIHd4qkrCdcAd+h
WEXPpqDaXcKf4RG/phiBw+lS/aLyFlAhZgy7H5MilBM/IAdaX21XAwfRR/WesMbt
O1YZINfhNFmfq1jQWHSBSZxsx0mDXbEVzIrbNxoTRcAFyQVbEdtLMUWVSBd1eYOh
96bxdcxymNlN0I/okdkDef2vlMMq9z463NknzNhXw91WubSdALDeLpZP9YYvYm1m
GlOiRLJ7/Ox4zhRYQezvjV7XsC45lKFMzuLbkbn3k9rE+U5BuXhgk+hGehFVXhMK
08fW+vVxfPnHGEbXr70+WnlrEM8oHuUkUxSkVAsZFGcKdnrTchINYsPXE/MnDnGo
VUdMNPTdD4gSE8Mx0pHuenKUfifgdVmwnZn6UpLSvOVIKidvVGmbPz5c1IMPyAcW
FxuoeyFGpQsvZ3FA0JTLxBxWV+nLvXtHrOGBdHDcCNXFs7i46dOuH1041bkCjLP9
E+f6+OSzzqfScr6w8Aq48uw5Dx7983FRQtA37m7pk1rfXEK5k3Aw0ayHlGpHqB0I
czHFAJ3G14RiSFIjctXzeMC+aAaBrEWuu/GQ8DrubUxwd9sHoiy607yOM4rJbqxf
imMeVqkM6tx1bgUXgrYDyMJVVVeW2sPDKZsmibbCJlsNf4MYHOHxOvZFMKs1E9gx
OMDtsBzLz2+RN2L4c8kmOBeOVIC/eraC1YHwvrGDIQR9JJKCGU0fGulTMkrQ61Jm
jcr090p+tSY4zZ2c7+W/zuAYINFrm6h7H6k0Bx0Fg9qjdWQwwq+Ai6MAL9brDJuB
hZ1uyRAtqAe0kRi32t+586h0RUIkvxXeTFYZjfQ52VZngtZDxujw8luS9LZBwNzf
lsa8U2IOmHTgKb94FFVspLF6dlE5Jd/tKJj0BC+d5PI4og3ONeskLq6veKGaCOfq
qzenfdZcnqgJ4Qa5N+bQtnF7ZOgLTzQkcwDA5DLkQy42U8chSY19cIgxzQ0k0ahr
cWUMU6xISGoa+RDzBvzmViuRamAjoPdoI7YKz2LLHIA+orHZzLvxJo5f+CleQoPY
26+Ft0z8nKGuha3fup4y4qVhlUYrCWRLL+6ZCRwBKo4uUtmq0/yqi7zb5uLfWoIT
UlD0uJg79eX90T8rVopKA3HPq9AtgIssiZ7GHK6IhWOeWqgx6sDsmJLxgfZA7z6g
3tvTbufAk5u4ZYYCHCczv979xJAbP6yKTYhfZb3R48bXbBCBBmAbZHS1/bllLJsT
SPuXT5XGp6zMzBGHolNHBzRGbtBrcbNXvSpVkTK+z5nDqLe6YiEyAyi74sUJCteA
Vi9R7sXCpaNeOxytldJdeTLgLRIAQuzsBeloH/iex1OSSdYpMrIhTpB0q2ibzLND
D0cj4uVleWV0oTRurdwqXJdNkI7h9rLLjLtUQFixzeI8wJAMXBeRDV7ugE+mxCYI
LbP44NQ3oCDY2knk6BTozjdy8AgPmuGm7kf9Xm866y+iH3x1LGiXscr1wBV7eMH5
XkTRcrQKSyMdMNoFDUOvBS4eFRydMAIzQ7HLyzB4ZtZuyE+e9jnm65NtGuWkFTXD
SOh9rE9IZ0P7pHasJa/jrMPTWBoPRBqmX+HpsZd1WZEtBg4+k3Zl7O2lt95uaj2Z
rn/4mIVWLT3coANiDbkn4XxBlZmpcs0oPFQqZMwr1iM5+4IOoZfxQI427k6iQrgD
6CxjA2fnmHhmLcMy1tyd+ciQYrk0F31uSBE89K4w+aSl6UrfdF0OgTC/Dd3oKYIM
KVlS6vde5x8NqSAbua//pRdMM15Su7r7mjCe7YjAGQHBEM0e2Ch7+jfB0icvpboe
Wnhg5TfqD8DkhB1aA6+Bh4RhhwcaaSZsSi+XtFWWPKA1wg+urqlUw0JlvMqfiO+q
3boGX0EDtplYA1981ELDrTguYHmmrFYBadSAx8SQ3kPc/3GL2KHJV03Ce99fx0un
1XQD3BoURmuNniMWle4ZQLMx/1UfO1tvnBajVe5KeOHlCvOsPvuM7VpLhGMiW7id
Iu8Mhi1feezQC9vaZZeTBTbBsvJ841rNWAgspI8nqsrOozZXQ1+qXQ681aP1B7BQ
Sk+X7lowWAjkrEqBEu0JFlu4WSAZ2Nkt7ju9Br6Q4fzQR2qxU9vm6P6EIkMUS5qI
sh3GlM7OGthe/9WfLqOvovE9/86dY6aCY7Phc0/LFUKz9QbSQOn9skkfaCvxLtsR
I/lJ7fV+Qa6+ekRxnyyxrsH7b236UCX9bBC4o+PzeVK5Q9zCHrcPgrJH5YPgo4Xq
NAbrlpovl1CYjjqPH5MF9TO2hBG2U1xjaegup2OEr9OZMXGq0go2rIp3pzAAr7Yr
QY808x5FhF5Rshn1G3Fe08YO8v/noHbjaQ+n/kXjOGFYmgkWNe174wmBDXqJi5Z7
IiQaeReWzLtU1ccQAcDnX1Slfyu7O76AKy4kpBhBmpy9Adn45eKxj6orUTPdw+rw
V2AKxw/iOBogN3XYf0eGt3INwH1EtBgrMZc7ppVkC7s5dkiHqZNODOkpRXoTXhfs
zKniQJ7gt9yIG0+a15MM3OD4SriF3flu8hm9SjAQeO6WxsVWBFR9dmpBDaXTrre5
+hlaYMelcx6nEcrUaSS+lCrT9+In6NYNZvrbloTclnSgqEhxIJFXA4CfM9gFrM7N
bdlldIkPYvb5qKYtDA5XHK1GVQT930xo94ci0YYsVfM5JMM5VBzH7ZeF2DIaUJnE
8UCq1SI1AZkAKdd7RwDZYIQEXjOvsHJi+BN295t3SUjBrhQidRP7uy303jvAYowC
8rdgO9mitG+o0w/gVAwJV+6+UPcsWpoSPBFboNroR0OCmIzLocqn5nfLwluBfYHu
oGoF7TWtyo4f4962WAleccnqyiE4w5cr5SLGQnOYct4K7DPOVlVxQxAgFi2HEIuX
/EkP+mBBCI0IzAsfTT+aoUxjbllTve0qo3Cnq/VtRiwIDLHlS4DUXnYvMyP4QbCU
fZXTITAebDjtbdbzSXOrjazFFQaW7YUgFpshDFnU0v2KNV4JvZ+RfSE4s97gLroi
JLWjJ1UNpTgVGqv5xx0uHPN/PyIaa1C5OJQcj4Y4SL1ly2Kb8n8CAhhcBXewIzWf
qK7hap3rD8dZRneDmibKMSMtrSIlAbhItJD3V37LxYaSC0jH7UQoIAuz28gD7HGi
xtD2b0crk5RQSTft9AsoB62qpGqrQMPtZMGpbMFvoHMSIzyWeMKp0IZOYTo1Tnxa
VTQxOdR2oIUZQAkpYr02ot+xQseiObqCqKrbHdNQN5xWSubc+wLkSeBXc8qgAAdE
JdYxiQAqAKR95Yj1Z/vz2NwRkdKaXw/YL104Pq2kjXg+Yiz6aDfxJ2hNLojOJYOc
0Ek5Sx4nygU5VXnVZKIfk8QmKi+ITJPC4GlX3gvTm08L2nre49n/0shiBeHqOjqX
79aGFUMnGppGF/B2tWLPQR9BVcnD6jXEx5hygMT3oYPmumwnXeSg6m04GODc3Ynn
6vvWEQw5gn20M8CRroJCyHILd0uhOFp9uMogg9dfctB70CGGzr7ViYJnAEUNYCSN
00tYH3f1dCxYEh/rTgEKGsaBoopwkb8Xqs8+c/e+DgPbeU+rWc4yodVT1R6Wk6G2
/MFTECAS1MczIMt1RmvPvX23PuHV/Mn/nGiA1zoLUGzNZ6HEG+gdXRrIWQRJ4L5/
bDnPqximsoDQJwXX44dZLu6YCl0dQoYAvZfJA8JdWUE2PyOmvafHrpxGsggMNR+j
fS66DY9ZQ+e125kkUNHgYQWqXEVgyW82MBUQ5KPPozexHeuD9WWd1gh6jxjBP4iK
ON4XycaC4v+sw7PJJ7tknbvA04URbDla9nPsAenpILjFzpIA2k4JNrmL3UUsgEBp
YC3PblqbsFxWsCx3xdSRXBSDP2z9cdX3Y6/RwIyIhvUll4iRk1ej7P+JEKmVyrWZ
6rdwT5KW2KTX1E5PaGG+EXFaMOWPwDBjZU2C8eS9HIPPXh/3adAEtSFAb9mRqx8k
`pragma protect end_protected
