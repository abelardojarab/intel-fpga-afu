// write_dc_fifo.v

// Generated using ACDS version 17.0 290

`timescale 1 ps / 1 ps
module write_dc_fifo (
		input  wire [109:0] data,    //  fifo_input.datain
		input  wire         wrreq,   //            .wrreq
		input  wire         rdreq,   //            .rdreq
		input  wire         wrclk,   //            .wrclk
		input  wire         rdclk,   //            .rdclk
		input  wire         aclr,    //            .aclr
		output wire [109:0] q,       // fifo_output.dataout
		output wire         rdempty, //            .rdempty
		output wire         wrfull   //            .wrfull
	);

	write_dc_fifo_fifo_170_bhnb7cq fifo_0 (
		.data    (data),    //  fifo_input.datain
		.wrreq   (wrreq),   //            .wrreq
		.rdreq   (rdreq),   //            .rdreq
		.wrclk   (wrclk),   //            .wrclk
		.rdclk   (rdclk),   //            .rdclk
		.aclr    (aclr),    //            .aclr
		.q       (q),       // fifo_output.dataout
		.rdempty (rdempty), //            .rdempty
		.wrfull  (wrfull)   //            .wrfull
	);

endmodule
