// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// Parse 4 word Ethernet MII stream.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_readmii4 #(
    parameter SIM_EMULATE = 1'b0,
    parameter SYNOPT_STRICT_SOP     = 0
)(
    input clk,
    input sclr,

    input keep_rx_crc,
    input cfg_preamble_det_on,
    input cfg_sfd_det_on,

    input [8:0] din_valid,
    input [255:0] din_d, // read left to right
    input [31:0] din_c, // read left to right

    output dout_valid,
    output [255:0] dout,
    output [255:0] next_dout,
    output [31:0] dout_ctl,
    output [3:0] dout_prb,  // preamble word
    output [3:0] dout_sop, // data word
    output [3:0] dout_eop,  // last data byte before FCS
    output [3:0] dout_eeop,  // packet terminated due to unexpected control character
    output reg [31:0] dout_last_byte, // last CRC byte location (i.e. 4th CRC byte) 
    output reg [31:0] dout_last_dbyte, // last data byte location before crc
    output [11:0] dout_mty // number of empty bytes in eop word 0..7
);

localparam WORDS = 4;

genvar i;

reg [3:0] din_is_data_r0, din_is_data_r1, din_is_data;
always @(posedge clk) begin
    if (din_valid[0]) begin
        din_is_data_r0 <= {!(|din_c[31:24]), !(|din_c[23:16]), !(|din_c[15:8]), !(|din_c[7:0])};
        din_is_data_r1 <= din_is_data_r0;
        din_is_data <= din_is_data_r1;
    end
end

/////////////////////////////////////////////////////////////////////
// if the leftmost byte is a 1fb then this is a preamble word,
// the next word is first data
// if any byte is a 1fd then the previous 4 are the FCS
/////////////////////////////////////////////////////////////////////

reg [WORDS*64-1:0] din_d_r0, din_d_r1, din_d_r2;
reg [31:0] din_c_r0, din_c_r1, din_c_r2;

always @(posedge clk) begin
    if (din_valid[1]) begin
	    din_d_r0 <= din_d;
	    din_c_r0 <= din_c;
    end
end
always @(posedge clk) begin
    if (din_valid[2]) begin
	    din_d_r1 <= din_d_r0;
	    din_c_r1 <= din_c_r0;
    end
end
always @(posedge clk) begin
    if (din_valid[3]) begin
	    din_d_r2 <= din_d_r1;
	    din_c_r2 <= din_c_r1;
    end
end

////////////////////////////////////////////////////////////////////
// 2nd layer comparators
////////////////////////////////////////////////////////////////////

// finish the 1fd, all positions
// JUST GATE FOR NOW - GATE WITH IN_PKT.  COULD CHANGE
// EQ BLOCK TO NOT ADD LEVEL OF LOGIC, BUT WOULD NEED MORE COMPARATORS 

reg [WORDS-1:0] match_1fb_raw, match_1fb_raw_r0, match_1fb_raw_r1;
reg [WORDS*8-1:0] match_1fd_raw, match_1fd_raw_r0, match_1fd_raw_r1;

generate
	for (i=0; i<WORDS*8; i=i+1) begin : lp1
        always @(posedge clk) begin
            if (din_valid[4]) begin
                match_1fd_raw_r0[i] <= din_c[i] && din_d[i*8+7:i*8]==8'hfd;
            end
        end
	end
endgenerate

generate
	for (i=0; i<WORDS; i=i+1) begin : lp2
        always @(posedge clk) begin
            if (din_valid[5]) begin
                match_1fb_raw_r0[i] <= din_c[i*8+7] && (din_d[i*64+63:i*64+56]==8'hfb);
            end
        end
	end
endgenerate

always @(posedge clk) begin
    if (din_valid[6]) begin
        match_1fd_raw_r1 <= match_1fd_raw_r0;
        match_1fd_raw <= match_1fd_raw_r1;
        match_1fb_raw_r1 <= match_1fb_raw_r0;
        match_1fb_raw <= match_1fb_raw_r1;
    end
end



wire [WORDS*8-1:0] match_1fd;

wire [3:0] in_pkt;
reg [3:0] in_pkt_r3, in_pkt_r4, in_pkt_r5;
wire [WORDS*8-1:0] in_pkt_stretched;
assign in_pkt_stretched = {{8{in_pkt[3]}}, {8{in_pkt[2]}}, {8{in_pkt[1]}}, {8{in_pkt[0]}}};
assign match_1fd = match_1fd_raw & in_pkt_stretched;

wire [3:0] match_term;
assign match_term[3] = |match_1fd_raw[31:24];
assign match_term[2] = |match_1fd_raw[23:16];
assign match_term[1] = |match_1fd_raw[15:8];
assign match_term[0] = |match_1fd_raw[7:0];

wire [3:0] gen_eeop_r2;
assign gen_eeop_r2 = in_pkt & ~din_is_data & ~match_term;

// finish the 1fb, starting positions (byte 7 of each word)
wire [WORDS-1:0] match_1fb;

// mask out if any of next 5 words is control

assign match_1fb[3] = match_1fb_raw[3] && (&din_is_data[2:0]) && (&din_is_data_r1[3:2]);
assign match_1fb[2] = match_1fb_raw[2] && (&din_is_data[1:0]) && (&din_is_data_r1[3:1]);
assign match_1fb[1] = match_1fb_raw[1] && (din_is_data[0]) && (&din_is_data_r1[3:0]);
assign match_1fb[0] = match_1fb_raw[0] && (&din_is_data_r1[3:0]) && (din_is_data_r0[3]);

// Implement in_packet indication; will
// go low if there is a control character inside the packet
// in_pkt_raw is the raw in-pkt signal that get set by start and cleared by any control.
// in_pkt is the real in-pkt signal that get set by filtered start and cleared by any control

wire [3:0] in_pkt_raw;
reg in_pkt3_raw_next;
wire [3:0] din_is_start_raw = match_1fb_raw;
always @(*) begin
   if (~in_pkt_raw[0] & din_is_start_raw[0]) begin
      in_pkt3_raw_next = 1'b1;
   end else if (in_pkt_raw[0] & ~din_is_data[0]) begin
      in_pkt3_raw_next = 1'b0;
   end else begin
      in_pkt3_raw_next = in_pkt_raw[0];
   end
end

reg in_pkt3_raw_reg;
always @(posedge clk) begin
   if (sclr) begin
      in_pkt3_raw_reg <= 1'b0;
   end else if (din_valid[6]) begin
      in_pkt3_raw_reg <= in_pkt3_raw_next;
   end
end
assign in_pkt_raw[3] = in_pkt3_raw_reg;

reg in_pkt2_raw_reg;
always @(*) begin
   if (~in_pkt_raw[3] & din_is_start_raw[3]) begin
      in_pkt2_raw_reg = 1'b1;
   end else if (in_pkt_raw[3] & ~din_is_data[3]) begin
      in_pkt2_raw_reg = 1'b0;
   end else begin
      in_pkt2_raw_reg = in_pkt_raw[3];
   end
end
assign in_pkt_raw[2] = in_pkt2_raw_reg;

reg in_pkt1_raw_reg;
always @(*) begin
   if (~in_pkt_raw[2] & din_is_start_raw[2]) begin
      in_pkt1_raw_reg = 1'b1;
   end else if (in_pkt_raw[2] & ~din_is_data[2]) begin
      in_pkt1_raw_reg = 1'b0;
   end else begin
      in_pkt1_raw_reg = in_pkt_raw[2];
   end
end
assign in_pkt_raw[1] = in_pkt1_raw_reg;

reg in_pkt0_raw_reg;
always @(*) begin
   if (~in_pkt_raw[1] & din_is_start_raw[1]) begin
      in_pkt0_raw_reg = 1'b1;
   end else if (in_pkt_raw[1] & ~din_is_data[1]) begin
      in_pkt0_raw_reg = 1'b0;
   end else begin
      in_pkt0_raw_reg = in_pkt_raw[1];
   end
end

assign in_pkt_raw[0] = in_pkt0_raw_reg;

//////////////////////////////////////////////////////////////////

reg in_pkt3_next;
wire [3:0] din_is_start = match_1fb;
always @(*) begin
   if (~in_pkt[0] & din_is_start[0]) begin
      in_pkt3_next = 1'b1;
   end else if (in_pkt[0] & ~din_is_data[0]) begin
      in_pkt3_next = 1'b0;
   end else begin
      in_pkt3_next = in_pkt[0];
   end
end

reg in_pkt3_reg;
always @(posedge clk) begin
   if (sclr) begin
      in_pkt3_reg <= 1'b0;
   end else if (din_valid[6]) begin
      in_pkt3_reg <= in_pkt3_next;
   end
end
assign in_pkt[3] = in_pkt3_reg;

reg in_pkt2_reg;
always @(*) begin
   if (~in_pkt[3] & din_is_start[3]) begin
      in_pkt2_reg = 1'b1;
   end else if (in_pkt[3] & ~din_is_data[3]) begin
      in_pkt2_reg = 1'b0;
   end else begin
      in_pkt2_reg = in_pkt[3];
   end
end
assign in_pkt[2] = in_pkt2_reg;

reg in_pkt1_reg;
always @(*) begin
   if (~in_pkt[2] & din_is_start[2]) begin
      in_pkt1_reg = 1'b1;
   end else if (in_pkt[2] & ~din_is_data[2]) begin
      in_pkt1_reg = 1'b0;
   end else begin
      in_pkt1_reg = in_pkt[2];
   end
end
assign in_pkt[1] = in_pkt1_reg;

reg in_pkt0_reg;
always @(*) begin
   if (~in_pkt[1] & din_is_start[1]) begin
      in_pkt0_reg = 1'b1;
   end else if (in_pkt[1] & ~din_is_data[1]) begin
      in_pkt0_reg = 1'b0;
   end else begin
      in_pkt0_reg = in_pkt[1];
   end
end

assign in_pkt[0] = in_pkt0_reg;

////////////////////////////////////////////////////////////////////
// checkpoint to eat invalids
//    need to see 1 cycle of future
////////////////////////////////////////////////////////////////////
reg [WORDS*64-1:0] din_d_r3 = {(WORDS*64){1'b0}};
reg [WORDS*8-1:0] din_c_r3 = {(WORDS*8){1'b0}};
reg [WORDS-1:0] match_1fb_r3 = {WORDS{1'b0}};
reg [WORDS*8-1:0] match_1fd_r3 = {(WORDS*8){1'b0}};
reg [WORDS-1:0] gen_eeop_r3 = {WORDS{1'b0}};

reg [3:0] din_is_data_r3;

always @(posedge clk) begin
    if (din_valid[7]) begin
        din_d_r3 <= din_d_r2;
        din_c_r3 <= din_c_r2;
        din_is_data_r3 <= din_is_data;
	    match_1fb_r3 <= match_1fb & ~in_pkt_raw;
        match_1fd_r3 <= match_1fd;
        gen_eeop_r3 <= gen_eeop_r2;
        in_pkt_r3 <= in_pkt;
    end
end

////////////////////////////////////////////////////////////////////
// reposition flags and start masking 
////////////////////////////////////////////////////////////////////

reg prev_1fb = 1'b0;
reg [WORDS-1:0] st = {WORDS{1'b0}};
reg [WORDS*8-1:0] last_dbyte = {(WORDS*8){1'b0}};
reg [WORDS*64-1:0] din_d_r4 = 0;
reg [WORDS*8-1:0] din_c_r4 = 0;

always @(posedge clk) begin
	din_d_r4 <= din_d_r3;
	din_c_r4 <= din_c_r3;
    in_pkt_r4 <= in_pkt_r3;
end

reg [31:0] last_byte;
reg [WORDS-1:0] preamble_sfd_err= 0;
reg [WORDS-1:0] preamble_sfd_err_r4 = {WORDS{1'b0}};
reg [WORDS-1:0] preamble_sfd_err_r5 = {WORDS{1'b0}};
wire [WORDS-1:0] strict_sfd_err_r5= SYNOPT_STRICT_SOP? preamble_sfd_err_r5 : {WORDS{1'b0}};
wire [WORDS-1:0] strict_sfd_err_r4= SYNOPT_STRICT_SOP? preamble_sfd_err_r4 : {WORDS{1'b0}};
wire [WORDS-1:0] strict_sfd_err_r3= SYNOPT_STRICT_SOP? preamble_sfd_err : {WORDS{1'b0}};

always @(posedge clk) begin
    if (sclr) begin
        st <= 0;
        last_dbyte <= 0;
        last_byte <= 0;
    end
    else begin
        // PCS won't generate more than 0x1fd in the same word ,
	    last_dbyte <= {match_1fd_r3[WORDS*8-1-5:0], match_1fd[WORDS*8-1:WORDS*8-1-4]};
	    last_byte <= {match_1fd_r3[WORDS*8-1-1:0],  match_1fd[WORDS*8-1]};
    end
end


reg din_valid_r4 = 1'b0;
reg [WORDS-1:0] match_1fb_r4 = {WORDS{1'b0}};
always @(posedge clk) begin
    din_valid_r4 <= din_valid[7];
    match_1fb_r4 <= match_1fb_r3;
end

////////////////////////////////////////////////////////////////////
// pack empty 
////////////////////////////////////////////////////////////////////

wire [WORDS-1:0] end_half0, end_half1;

wire [31:0] last_b = keep_rx_crc ? last_byte : last_dbyte;
generate
	for (i=0; i<WORDS; i=i+1) begin : lp3
        alt_e100s10_ohbin8 ob0 (
            .clk(clk),
            .din(last_b[(i+1)*8-1:i*8]),
            .dout(dout_mty[(i+1)*3-1:i*3])
        );
        defparam ob0 .SIM_EMULATE = SIM_EMULATE;

        alt_e100s10_or4t1 c0 (
            .clk(clk),
            .din(last_b[i*8+3:i*8]),
            .dout(end_half0[i])
        );
        defparam c0 .SIM_EMULATE = SIM_EMULATE;

        alt_e100s10_or4t1 c1 (
            .clk(clk),
            .din(last_b[i*8+7:i*8+4]),
            .dout(end_half1[i])
        );
        defparam c1 .SIM_EMULATE = SIM_EMULATE;

	end
endgenerate

reg din_valid_r5 = 1'b0;
reg [WORDS-1:0] match_1fb_r5 = {WORDS{1'b0}};
reg [WORDS-1:0] st_r5 = {WORDS{1'b0}};
reg [WORDS*64-1:0] din_d_r5 = 0;
reg [WORDS*8-1:0] din_c_r5 = 0;
reg [3:0] gen_eeop_r4;
wire [31:0] eeop_last_dbyte = {2'b0, gen_eeop_r4[3], 5'b0, 2'b0, gen_eeop_r4[2], 5'b0, 2'b0, gen_eeop_r4[1], 5'b0, 2'b0, gen_eeop_r4[0], 5'b0};
wire [31:0] eeop_last_byte =  {6'b0, gen_eeop_r4[3], 1'b0, 6'b0, gen_eeop_r4[2], 1'b0, 6'b0, gen_eeop_r4[1], 1'b0, 6'b0, gen_eeop_r4[0], 1'b0};

always @(posedge clk) begin
    din_d_r5 <= din_d_r4;
    din_c_r5 <= din_c_r4;
    din_valid_r5 <= din_valid_r4;
    in_pkt_r5 <= in_pkt_r4;
    match_1fb_r5 <= match_1fb_r4 & ~strict_sfd_err_r4 & ~gen_eeop_r4;
	if (din_valid_r4) prev_1fb <= match_1fb_r4[0];
	st_r5 <= ({prev_1fb & ~strict_sfd_err_r5[0], ~strict_sfd_err_r4[WORDS-1:1] & match_1fb_r4[WORDS-1:1]}) & ~gen_eeop_r4;
    dout_last_byte  <= |gen_eeop_r4 ? eeop_last_byte  : last_byte; 
    dout_last_dbyte <= |gen_eeop_r4 ? eeop_last_dbyte : last_dbyte;
end

reg [3:0] gen_eeop_r5;
always @(posedge clk) begin
   // Do not shift EEOP back; let it come out right away
   // Gate gen_eeop_r5 with st so you do not get SOP and EOP at the
   // same time for malformed packets
   gen_eeop_r4 <= gen_eeop_r3;
   gen_eeop_r5 <= gen_eeop_r4 & ~st;
end

assign dout_valid = din_valid_r5;
assign next_dout = din_d_r4;
assign dout = din_d_r5;
assign dout_ctl = din_c_r5;
assign dout_sop = st_r5;
assign dout_prb = match_1fb_r5;
assign dout_eop = in_pkt_r5 & (end_half0 | end_half1 | gen_eeop_r5);  // word with last data byte before FCS
assign dout_eeop = gen_eeop_r5;

//---------------------------------------------------------------------------------------------------------------------------------------------------   
// UNH compliance - START, Premable, SFD checking
//---------------------------------------------------------------------------------------------------------------------------------------------------      
//
// SYNOPT_STRICT_SOP = 0, Default behavior: only check START. If START check fails, no SOP generated and EOP will be handled by downstream logic.       
// SYNOPT_STRICT_SOP = 1, This is the new added features built on top of Default behavior.
//    0. START is always checked. If START check fails, no SOP generated and EOP will be handled by downstream logic.    
//    1. Check based on MAC Rx CSR configuration 0x50A[4:3] = {cfg_preamble_det_on, cfg_sfd_det_on }
//    2. Please note premable here means 8'b1010_1010(per spec). We don't check against users data in premable location when in Premable pass through mode.   
//
//---------------------------------------------------------------------------------------------------------------------------------------------------   
//
//     +----------------------+----------------------+-------------------+--------------------+------------------------+-------------------------------+
//     |  START Check         | SYNOPT_STRIC_SOP     |cfg_preamble_det_on|   cfg_sfd_det_on   |   What to be checked   | Behavior when check fail.     |
//     |                      |                      |                   |                    | other than START ?     |                               |
//     |                      |                      |                   |                    |                        |                               |
//     +----------------------+----------------------+-------------------+--------------------+------------------------+-------------------------------+
//     |      FAIL            |     Don't care       |     Don't Care    |    Don't care      |    Don't care          |  Default behavior.            |
//     |                      |                      |                   |                    |                        |  Ceasing SOP.                 |
//     |                      |                      |                   |                    |                        |  EOP will be handled by       |
//     |                      |                      |                   |                    |                        |  downstream logic.            |
//     +----------------------+----------------------+-------------------+--------------------+------------------------+-------------------------------+
//     |      PASS            | SYNOPT_STRIC_SOP = 0 |                   |                    |    Start               |  Pass SOP EOP accordlingly    |
//     |                      |                      |     Don't care    |    Dont' care      |                        |                               |
//     +----------------------+----------------------+-------------------+--------------------+------------------------+-------------------------------+
//     |      PASS            | SYNOPT_STRIC_SOP = 1 |                   |                    |    Start               |  Pass SOP EOP accordlingly    |
//     |                      |                      |       1'b0        |       1'b0         |                        |                               |
//     +                      +                      +-------------------+--------------------+------------------------+-------------------------------+
//     |                      |                      |                   |                    |    Start+SFD           |  Only pass good packets.      |
//     |                      |                      |       1'b0        |       1'b1         |                        |  Drop failed packets by       |
//     +                      +                      +-------------------+--------------------+------------------------+  ceasing SOP and EOP          +
//     |                      |                      |                   |                    |    Start+PREAMBLE      |                               |
//     |                      |                      |       1'b1        |       1'b0         |                        |                               |
//     +                      +                      +-------------------+--------------------+------------------------+                               +
//     |                      |                      |                   |                    |    Start+PREAMBLE+SFD  |                               |
//     |                      |                      |       1'b1        |       1'b1         |                        |                               |
//     +----------------------+----------------------+-------------------+--------------------+------------------------+-------------------------------+

//wire [WORDS-1:0] match_SFD_pre;
reg [WORDS-1:0] match_SFD_pre_r0, match_SFD_pre_r1, match_SFD_pre;
reg [WORDS-1:0] match_SFD;
reg [WORDS-1:0] match_preamble_r3;
reg [WORDS-1:0] p_preamble_high, p_preamble_high_r0;
reg [WORDS-1:0] p_preamble_low, p_preamble_low_r0;
reg [WORDS-1:0] match_preamble_r1;
reg [WORDS-1:0] match_preamble_r2;
localparam SFD      = 8'hd5;
localparam PREAMBLE = 8'h55; 

generate

if (SYNOPT_STRICT_SOP) begin: gen_strict_sop_chk 

	for (i=0; i<WORDS; i=i+1) begin : lp4

     always @(posedge clk) begin
         if (din_valid[8]) begin
             match_SFD_pre_r0[i] <= (din_c[i*8]==1'b0) && (din_d[i*64+7:i*64]==8'hd5);
             match_SFD_pre_r1[i] <= match_SFD_pre_r0[i];
             match_SFD_pre[i]   <= match_SFD_pre_r1[i];
             match_SFD[i]       <= match_SFD_pre[i];
         end
     end

      always @(posedge clk) begin
          if (din_valid[8]) begin
             p_preamble_high_r0[i] <= (~|din_c[ i*8+6: i*8+4]) & (din_d[ i*64+55:  i*64+32] == {3{PREAMBLE}}); 
             p_preamble_low_r0[i] <= (~|din_c[ i*8+3: i*8+1]) & (din_d[ i*64+31:  i*64+8] == {3{PREAMBLE}}); 
             match_preamble_r1[i] <= p_preamble_high_r0[i] && p_preamble_low_r0[i];
             match_preamble_r2[i] <= match_preamble_r1[i];
    	     match_preamble_r3[i] <= match_preamble_r2[i] ;
         end
     end

	
        always @(*) begin
            case({cfg_preamble_det_on,cfg_sfd_det_on})
                2'b00: begin //check START and SFD
                        preamble_sfd_err[i] = 0;                              
                        end                   
               2'b01: begin //check START and SFD
                        preamble_sfd_err[i] = match_1fb_r3[i] & ~match_SFD[i];                              
                        end
               2'b10: begin //check START and PREAMBLE
                        preamble_sfd_err[i] = match_1fb_r3[i] & ~match_preamble_r3[i];                              
                      end         
               2'b11: begin //check START, PREAMBLE and SFD
                        preamble_sfd_err[i] = match_1fb_r3[i] & ~(match_preamble_r3[i] & match_SFD[i]);                              
                      end                     
            endcase
        end   	
    end	

    always @(posedge clk) begin
    if (din_valid[8]) 
        preamble_sfd_err_r4 <= preamble_sfd_err;
    end

    always @(posedge clk) begin
    if (din_valid_r4) 
        preamble_sfd_err_r5 <= preamble_sfd_err_r4;
    end

end
endgenerate

endmodule

