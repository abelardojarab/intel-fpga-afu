// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// 15 bit val == const(7ffb) equality comparator.  Latency 2.
// 17 bit val == const(13fff) equality comparator.  Latency 2.
// Generated by one of Gregg's toys.   Share And Enjoy.

// 17'h13ffe = 'd81918
// 17'h13fff = 'd81919
module alt_e100s10_eqc17h0007ft2 #( 
    parameter SIM_EMULATE = 1'b0
) (
    input clk,
    input [16:0] din,
    output dout
);

wire [3:0] leaf;

alt_e100s10_eqc4hft1 cmp0 (
    .clk(clk),
    .din(din[3:0]),
    .dout(leaf[0])
);
defparam cmp0 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_eqc5h07t1 cmp1 (
    .clk(clk),
    .din(din[8:4]),
    .dout(leaf[1])
);
defparam cmp1 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_eqc6h00t1 cmp2 (
    .clk(clk),
    .din(din[14:9]),
    .dout(leaf[2])
);
defparam cmp2 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_eqc6h00t1 cmp3 (
    .clk(clk),
    .din({4'b0000,din[16:15]}),
    .dout(leaf[3])
);
defparam cmp3 .SIM_EMULATE = SIM_EMULATE;


alt_e100s10_and4t1 c3 (
    .clk(clk),
    .din(leaf),
    .dout(dout)
);
defparam c3 .SIM_EMULATE = SIM_EMULATE;

endmodule

