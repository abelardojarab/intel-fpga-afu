
module pll (
	locked,
	outclk_0,
	outclk_1,
	refclk,
	rst);	

	output		locked;
	output		outclk_0;
	output		outclk_1;
	input		refclk;
	input		rst;
endmodule
