`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Mo7zCaZmS2Nk9OYA1PKBeHL4WbDTS3kf3T7nvZFKKTOdILiwG3TUqZIvIvl99D/2
v/EW5F0vj/I76kcjle7y6+t64ns6GMB4+91idzvroy9wuKpBoR81T8ZaDaNqunM1
aygO8XoDhD8emXdCbCeS2YHpZEMk+PUoMzcAYyN9T2k=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6288), data_block
wwKP/RwovevPmLDQgJ4C5LQQ+cP/SMeYaIMhAty0O15GTKCOdqB/jiKeZrXQlaPV
uZtmSSQJ+MEvgFsHQzLWtaLV+YsuBQs7lmnuIGJoKn3gs9o6ijPMBIz0JKeiN0rH
aspAMzQCuqdv79oYxtAHs0Dl3DkO70lQAiNxG6nZSOEXOjKguv8mIuZB0djFXjE1
32mK2HDhJzjSzL9dXxYN9aaRyt5D8Wrh41dS0ia1PGnmzBYJN6VlZAM9YoaD1wYS
zyCmuA6hA8gDjw7FyJLwkE14aeNMnvrgkZmKNSUNN7R3i7FZCUrI20lLMLc9uIV/
eX+IB+q2Kmsy9qu+SmtXGb355x/Icmfv/Kk88Wcs7b1WB/zh/fUs4BQQOlSkhCiS
3rU4JThaauZi9d1M/J22V5MI+VcMxBeqG+CAHGGpg668H51I2ZyHhLHUWdcN0iQb
FJpOSmVHFV3TGJnW/wSLUwvpMLBzQt8o+Jc2ovQzRQQ1CxSPIm+a7IrHyFTb5I1b
Y7kWGqpFvJ4SvaS1+lwXBc2auiHJnsOxKHCa7fE4n+oYvzsULT7KAv9Mo5ZLP1F9
sUrPBcv2kkMwhUe7leGw6N7oe1G8/pM5qz0F4RMweNSoD/BsUOyAadUAv8HI87yW
g24IEkDhxe2udfCSLiNPZ+Tw1UeuEptrK0LCQJNAh/cSgaQmMXAsix/qnbmqhp2v
RJSOidyz7nhqauIDMoJ4TjJH7K70BzD5K3f6n82mKbE7+SRyNloNf45ajXSoc1yU
BR6Yaafha6pNlRJ7NawiOfn6Paw9cigOPbJdMT3f1JpkAHpd1usUjOtvh9JDuTEQ
DMfY9xV64xi1raloCfhY6DVEFrW9bxK5gbZFItlV6WbeMGnnkMjRSbM6YTggvHcU
RFg50OZvyZ8UTwNnfzGf4pJSAcs2IyXmhn4di0+Gl2MpvVkOk1UCqMdQVLaWQYyJ
hA0T5rPP/IoIhzZdVmdSeV4MrmAuDRaXUNtktdKL4qwPQnKUy+4bnwXevspRV3HC
fOzaHsUVzvIIQMeJWbSqoia3eA4SdNSLLzsTFH8Bt2FgDR8hxhn244IdvDkjrrsr
yIPImwjwxTWXV+VDzmetNGwyV4ywRSCuV4gPxzEyU3r8GdVJ17qlZF21KPhMjfWg
phBloCON2rDgmWcRlNugyFEU6bjwRrOGvkYVns93FL1Uo+Fbz7ztwbwPZ6Tj4+6T
ppAuM9MQuTy1mTKkSp5WD1D2bECGJVwpr5Fy06uHi/HgnAQWGsHAbdcIsHenpjqw
1FN+UhZr+s2MkfJDJYW+GBAEd2mZ6GvQj8tcs3fjptzgzt0IrYYJHt4E2KdA5Uo+
DeGWELSgnGOwb07La9h31iWodIEENM00MZLyK3EBDnHwj7OH51xTWNwzUtS6DBDB
30Ity4sn11Ti1LB3frQKUqh7LE8v+q1F7aMHk9h4+LldWY2l61lB8WLwmxIyTSa4
Ll+ogUFm4/q0tHlZiy7BNg9hEe14hF+EmEZrXx9OKw6XvSO7ir1Nfw110ilbU9Uy
Iy0UYGxHZnkk4GjuBpWVEf2rzBLNsxy5JgP2xqNJ/PuiYF//3QJh5faKAYxBWYEE
uZCsaIoTbmMEIMk+9TjWy8krjzef1k7wF1XQ48/eU+Y6300CCLAQiBabQanLyGC0
eMu9aMy8B1Ew0KKQYJlQTa7rUUpJLXHL6+aU1wA6KvubXRoBdvtRQokoOvNfNfYF
Gw0uaPm6Znx6U5vqypgBDEJOU8oNLd4NDtGuQc+2JSEkcnTc9VHn6Wk0m2DTf/dx
HFuGeatHPsB0LS/6uwLax+L1+DjMFXzYRlvQlyuKKncQkScaVHtuD5A7M6aEsmr9
0c6iVhnS5paF+N++jPp13Q7fl5e21d3ConPb49+7houje8KwrlwT+XMnv4fdKskE
tcs6yb2ganVGt6rYs44jbDb2hk624emTK8z1mTjG5JBsNVnpeL0eOG0azVYUpAef
Tj9yRkCfYBNAJQU8wW3Ifqs4p9xhsWYFIYjRnKqhu/+nkn8cTera3p03wPhOQvtw
HtAzO2VBy0OQ7Or7ai1y+JsJF69ssO70QOPCUH+l82rbRRpTsjfVdzxo/vXx9vsF
R+RcT3gMDQetGylpOxkTEpeZ+JF2xUEpAvBiPhQFS49uN+Czh2oYtbRUWiffuABA
6/ARqNTcktihsSrxWZLsifZg5Z1zk3GPIVGvMt55jsO0YTGJ1+d1cOr+Lz76C0UJ
yFLguiVmUm9NorBZpd8gEw9JipgRYAlGR+qypVEeVF78Ace3cjG44jSHYB31A0bJ
p+YnjjSfOqK78Xpos55hgu6/ziIjlSAUftO9B/36ubEMjLPpXx+q9wWWTEHgYQHW
AhYCf+LdaxyOmt9VMVCt1bJfzvT7VhKsPD5GLOrxYUxW5ycTuVCJN7nG/8bCUZfX
ApIOqiVgwhAmyS3bCtL6NYnl5h+uoUqvj5PPlAAUmGm0cE7QywUKShbBvRbj+oZ3
I3EBDtNh8JhaCaWDk6XeZsm/4VpJFtFCBAnqlNH2P6T/PKBG/QCsm3jPGeodGxfp
t1jEd+Qz1uae0vEFhy1XNqMxXQ7l2DoQ3GAPK21WcHMO6VD7e4UvKvVSGAFivkvf
6fE7Yqo4Fj5jmMekTLJy+vXwwxu4LfMhwsAEBHaRul88g6l0oWVTO8cdYMTFjaGP
bi1Owx9zu3OYo/UUfoxPCBk+zHG7kkpe9Ewla17y4MYbjGMEaVBGdWk91/xRPZWL
I8iEc+X8mH/j9s9JS3xY6oENuy1lCcLv46LFsR80QX1dQeKeL32IkzjPiObLyxeL
g5DPMy9Dd+ggCQ/6iBRoZkUF/GeAvUJiiIrJnS719nKxIvsYSZWWq2ds9Fx0IqSW
2sKwnNDkqM2eoLNKPOj0P1ArD7XI8dSLk7CylY85g821ohZVkX6tAoL6Rp01GOS5
bexO/dEE0dBTgSWZWF3W/ELl1SznMPjPlLZvVApAfcg0PTgCtiZVDTNGZ9m8VyKs
37X6PoBnHf6GsnAQ0tCFbxkQz8L6jZPFk7pWe0d/FFLfdv751QsTwXI7mKIjdUVD
ulDMR1N70Ggr7yG+ga1dVqmF/QGpb8BGAlHozMJdged0y1wTcq4Hjx9+SHQltIw3
qOp3aSz98mwFJPKqdYpy02vHSbHW30ZXP0Cm9QoA9xvz0e932tq6nN4c+/IHHJ1S
eWKEabtEZGrpsi4s5nWZ94v38VUTSuMIOAR1+qW97rh9x+D1DPiTqxpgpmKRbdHv
YIfGNBOez/yyq/ZWTUtM1mpPjc9WwhLKEYPJaY/npMlst0Se3pv9rdIIISJGTq5q
a6lSYEfH809kHqisHlIoZlo6bXZlr/qDs1vR2cQoedJ8k5nwsSkKcTAiPoFYMpNv
lN7wQlMbStAy41byMfaAoBKiCUgo8fPc6AJzxU1oi73YaNwJdB8hl0kcND92QbId
YgPy/vg8bwA1KoK1JgLGO39zBUkt6uMgs0FO5R9n0cqBz+XGKTEebJeQ1UPR1G9u
oKbjJ/3xz/krkG/VupoyrixblFdxrHMkE4lt5G/EpQ1UnxA8Up3uWK3byUzEhaej
5P8jI+Ab9dK7a4vFwDSM8J9jwBii2y4SU1RWDFoOHPq51TUOg5aV78reEjxtvuWs
apkxbJSSsA46lT+q9oxPoYIVnuSUno53MJ6JWPKWHHPLutd8xxaj8xru8eRpHR46
7+GjFWjy8OAHDc0n2MVxj1HSqL/6JdcgbgQRvD4PuIpDfGcaBRtdgEyo0+ellINM
x21XWGjeWEQGfZBNeDp+e9MJSkZ7UQxBLU7c4Q5XWauHZjN9obQtBuZv+wuWEwUv
Oiazb1T2Zmjzdn4SfSCD6kqIooklJB5orEAX/ntF0zG5oYSlNCdv4C29UV/YUtfw
ilk6OSTuYTTWamHyY2eiheTqb6mr1t7OxydP3nY+lYTiMYQBWk6NDTGEj1h37GGq
LUBsHXV18h8thv1Pk9CNw3GfrI5BWWoAravxQdTLTf50+2gTHJ7v8N/mH+Ho9JWp
6eAUQcTRbDXnoSCVMZDysEd+aiuLEUfjgIXaVZCjaNI2I0fagYkKLTDo5fl49v0o
QtAau7Dq7xuVO02nVTb47WlHWq31BlwzeimvOXQt6Pq6x8whX7i5cM6gMsD5li2L
nHZUTWxDqrm8sB/+RcREwcd63awv3elKqaLQWil+ps3sVkJvh5/ao4q6ho5OfW50
IuFThxszn3a9BCa5Msx43WoWf3JF09Qxgq76f7ZVH5EY8o/FGHLnKxFRpfpWwDZK
zdzFlhHGm+ptffsmljAAZ3r09wW+uzQksKQVcFPlLJOPJkRB0LYKhz/L/Qs+G1nP
PqaSh6ArfgacrTakkZwrc/DeXizt7lbMqN9r0d9elwp06cxuHQUqYIfMTzEjIBBd
HDJlQ6Wkeoh6XQwNuT4XOADA0M8TQtsAnQ1qUUuNWkreLdziMNELOBTNdG3nuGZF
USkcX0GQovuHCZlT1tn8u5PTSQ3XMYa7HWRRXuziFOSPl10ja72RG4bZ1SL8iQKf
yASjD+xJffs4toQSJ3WjNVChSJcK3lkWQ/UXKaeLUSrulBJTWm4/FGyC/Assb5pD
t4AQI5+pTE7QmVBhJNAvFin+tzV4rUj6c2x0Euuy/RbGyogaTWC1eYn6mKWZWzEj
51y2EU12I8rBZuB8bHWTbpGVoGvDxnHphbOy92YUMYeaxumjXHbSRFtgUrzqL1pR
zKkWeKw4I1EYEBP0LLAq9ueseEQoSYcY8Y1Z3r8i2VTouXwVwymuEGeONVIq9DEI
s4eTn/XguJuKzm5I6fE04fWisIcbvBeRiMzMC33SKFwUB/jYYMSPWC3U5o19/gzR
Yxu3LWD7h9PcbZGX7V5ghew6FJpkbn0KwYwHW/jsMC8cjAVMgLcsvpGY1kX0kaLh
Ez4NnVTvQd4s/xe9AZrYrEUi557PAJ1ysrAccbkGbpLZeQaXb3tB/wlBS9MEaUTj
Oe+4LFzhLST/2ISXk3iyzqHemLNZKUtS3bxrirTLyL3Z6oOHUuHp4G4/AYsHgPM4
JXjgBBWtkJ7t0pVIZO2ICgpGdPTr2Bk0yYnWRic9jeu2MDoP0Dwldp73yQzGcEZJ
beBLRKUP9qIGRQHSKpYpgQhpRGA3d4riu8iEinpeukgW9c8Fe/lLeoWMezMKsjAl
ReWdho7gK1zvk7P7IZA2/iR5S/DovWyeAoDj6mbQBuRz3UubkO6TiO8oh5PTH8la
HhQng43FWkABQCd7qTHpH0dSdiDKfeypKwBr0cAAIFF8+qWWJxJUa5jrgnlQXiHh
d+CbV9gk31IjEoKs8BlLTI37vZgBEqsqMLqxgZojLgxVe3UbHzZ5KRACip6LJ0fX
Sm9oIyxTwbTHO9pAsFFPFtpzhKybDbZFmFwcWnHs7p6VtYLToRujLzxmQ5m+/W0J
7O/p6hkrQsuB4QS8yNf4OrzJO/GEfHUqVIuCWNxHRBMV+M/g/kRfYA1/S2so6dpP
BN8iQ4QOi1mdecqEuZKpP+6sYPsrl2/elqAIYxcog6ZkzIukb2zgVBhhRajVi05d
XG42B3oIbAzWX0+qlzJTYTDUurKYJ94ZYqns9He3p7UABCTda80RvTjJvRdncBAA
8J0lYNqSTCQz0TUr4yiPORx+FJkB1NYiZJxTD9zZzXROfyRJ78DoneluaTNZ/P6t
pbJo8uxMQ6Z1PpFv61rw4ryBtU8ba5yf0QtiJw1JhLSGJPMdCyY0jHmOSKj3EN5E
lZOHS1ka5q46L18RiaRkj7iFy5B/L0kVxm4KkJAjxLVoc9jjH+1VWXRSUHCIX0xE
nGnfmHv916PfoOaMyMv/NmqLGYevuUqE9yZQrbsbSPf05sFE2nJlQQfe//Z4z2a6
THEVwvfK+1kDJGDlFocNhHe8X9LBHyO9qoUZI5z7aPhmTOrgX1rWNhvC2O0a+YnZ
1cPJsktTUWaITqzsuyTrEBGvR2Lvjz7lBgEiNIf2CjD91bYRDlNoABz8h4DefNoC
5LohsBJB1TZrTWq5uPFl9kdxPDbsYbrGE3iS+sAc0XHtnbmV7obFRCiHg5hAqIMP
Y525AyujVNvFgfya/ig11ldFawdNDI5KHsuFkj/z7oUZy2URcPvISyta3pCuOs3C
HYQX9+KH8ypd7UyWHKJDV3auWv3EmAeBYOjVAkJgX1vZj2YfTH3SewwYfQ352WvB
VGSnX8vxZU0FlZhvTFbY3uiJ8QoXeM3hSqfCsHCNptDZ+ShNi+6wl/EuW3UkWQnU
NZKWiBIExHmcyRDLeGsesOIpuyVQIwxcjj8xL18IrFxLbCjjxP/Q22pnwjgHHMXD
V1i8aj/ImIUaZfj9IBUs0+z5aA3k1EigKEZdfWn7W8sWDDLv3UNxziQh9ipEkTpC
TDMrCgC/kKMD0FYD/9FOBEl+PsawDh27Dg8NDiBJbvi9NQ0OXe4w1jqz3bUR0ls+
q8IbyYRYEM3H941tpIjNt1CaN3pznp78Ywzf+EoC7+XC0mth+w6mPCdxCTrrMGNt
NIVaM6SNNrqE1wE5nIAQG1NHN0xxV8w65GS8fOGK5iIJHsjyxCcnYovPAbM+5Qfo
MH9mWG+VONT5cWBvdgs5sagzyRfkPYVTvQN8U+sQwSjhzKQCo0U1PqqROW8KBNVk
+Yj0UsoDuUa823IXv3hwHA4r399ccAtL/SrNFkfkGg7q8nd5ljXW6iwKqCqpeNTI
HHt2LJ+hojQAb1dEHA58ABmdGR+5+khCrLdVEkvmfWuMhb6B6TJW2HAuwUzQgh9j
66CzZsYHTrU6SEpb34GJNk15d1GkaG3SKLb0MC9+IBt6LLMIqM2isdxSoGrQGk8y
nUtuhJcZDoeL6u28iwQEXaQY4NqzCr9xuhEv3SYEKdv42ncqcoh9sQYKNRxIx1r5
QeKD9S12xeHMQWYaF+w8zqMX5YE8HJv3WqsA3aSwZaL5uuF+6Bp7o50Nzb04LsZm
uLotgw2qNiiDsaFkCIi6FtS5cYWHJI/jRohH6N8Wur6mEwL0dg/h8uIfFP5RL9Ir
Wrw3hSyjCYmGYEjWxFJxznMaFBkouK6HYzAJoGst1soPaby60gPXkmJscL6TUuBK
KubuFID3IVygVMdG0xYyOCo9bgP6KnZ8uOWUJEL078FDp7KEcpqI1RAQESRNE9/B
HqNoWeQP6eKdwx2TymduswIfqmM+Ur1pCDBuUx2NIKabKKXZzJ/ZThW1ogaCkRwU
W5CsXlKy5u+6SAb9IYP5/bD2FT+6ALaxhzmwuyqWPCUWKy7PYb8j33+qbHbx3n3P
18arpcgJyefFKWGeu+xjtaj+9gs7ciWdR3VlffEktNYWhnSTFzy2k/GX7BTE7qdN
qqXcIxCiXRon5UPk9suAddonqcdsrakyw2ceOK+YHluGfJyhzfpmfo0RW9BiMBPo
Yht+YX5fN6wn23iXzQ9xsVG81yeIy2gK4dOmPgv7bcfzOfE7lmv3pyYYeY7Rl1ec
hUrKQl1chZ3SIw/9EOET6otrYpEZ7Xr6ClOMNy/8yhcilAaP0TONGJr3mf7Le7ax
AwVNzTxoo0psQZA24jB6w3Kw10Qfbl6OTVyBfO70dI4c2A+da1R/SV5r6vhOanEc
9XZME40KmZ445WvqKmLbXpWt0dajHewySQY7AaSfIO7Aa3mnJUJJJN0nqY+8SACY
WUkCrKZjG3nJEoRjWslA3sOZka4n40i+qdB+ZVvEBQJTecgRT22WoX6HlQqvtCwP
s/fXNwc7CHgJyj5MihufJokXu3Co2wuCEp8wqeDRr1Ywm5/NQT8Qy4E651FqNygT
8MVLA3My718qO7N4GJKna4NUFZZF0cmK3gKyu3hAa3EkiCNJnmkVtCFH/7jEHQkf
jo11NcUMEBb55/03E2XQKRsrCki7+JhIFOdi1P8FrZy/NLLUrihMcQ/fFs8tbg/Q
9er4rajAjAXNbNTSelAG0iB3kOT0j9OuV7wGTGf836nzET16417jtsc0fr2b6zOz
/3Zsd2drWOatqMX0wwOTTo2KVBybK+0HTEuooR/69FeBbrNpYjO8JGy8g+k+OoNR
+SOsIOWOjVGH30x3Kk7YDgd8J3nLdM0uTjMYAzdZmaymMJYabyHl+4uzHnB3gP3V
hEOCvTw9ng61OG5WFWxBIc2hMdvcUPAmA05qGHQtDhGNZxwrwVFYa69R+7Ie3sRH
n55YYAaAGhwRHauspPbpHsRmL0A2bqblSs2n9O8734ge7Bz7tSab9QUmtviafdPA
o6In6nymswM+fUV/mfFKHqD5sorOr991SVEEVcGD8Z+Bcp2BHfhUmrV2nS1+Ppj2
dpvSzLkcfAJQRLTtyyXZqleIZS4nyANn7VzWbZWGkN5EUMhmb3EMZ+njftV+MDwJ
`pragma protect end_protected
