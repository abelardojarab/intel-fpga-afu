// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// Opposite (A==~B) compare of two 33 bit words.  Latency 3.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_opp33t3 #(
    parameter SIM_EMULATE = 1'b0
) (
    input clk,
    input [32:0] dina,
    input [32:0] dinb,
    output dout
);

wire [10:0] leaf;

alt_e100s10_opp3t1 op0 (
    .clk(clk),
    .dina(dina[2:0]),
    .dinb(dinb[2:0]),
    .dout(leaf[0])
);

defparam op0 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_opp3t1 op1 (
    .clk(clk),
    .dina(dina[5:3]),
    .dinb(dinb[5:3]),
    .dout(leaf[1])
);

defparam op1 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_opp3t1 op2 (
    .clk(clk),
    .dina(dina[8:6]),
    .dinb(dinb[8:6]),
    .dout(leaf[2])
);

defparam op2 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_opp3t1 op3 (
    .clk(clk),
    .dina(dina[11:9]),
    .dinb(dinb[11:9]),
    .dout(leaf[3])
);

defparam op3 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_opp3t1 op4 (
    .clk(clk),
    .dina(dina[14:12]),
    .dinb(dinb[14:12]),
    .dout(leaf[4])
);

defparam op4 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_opp3t1 op5 (
    .clk(clk),
    .dina(dina[17:15]),
    .dinb(dinb[17:15]),
    .dout(leaf[5])
);

defparam op5 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_opp3t1 op6 (
    .clk(clk),
    .dina(dina[20:18]),
    .dinb(dinb[20:18]),
    .dout(leaf[6])
);

defparam op6 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_opp3t1 op7 (
    .clk(clk),
    .dina(dina[23:21]),
    .dinb(dinb[23:21]),
    .dout(leaf[7])
);

defparam op7 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_opp3t1 op8 (
    .clk(clk),
    .dina(dina[26:24]),
    .dinb(dinb[26:24]),
    .dout(leaf[8])
);

defparam op8 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_opp3t1 op9 (
    .clk(clk),
    .dina(dina[29:27]),
    .dinb(dinb[29:27]),
    .dout(leaf[9])
);

defparam op9 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_opp3t1 op10 (
    .clk(clk),
    .dina(dina[32:30]),
    .dinb(dinb[32:30]),
    .dout(leaf[10])
);

defparam op10 .SIM_EMULATE = SIM_EMULATE;

alt_e100s10_and11t2 c11 (
    .clk(clk),
    .din(leaf),
    .dout(dout)
);
defparam c11 .SIM_EMULATE = SIM_EMULATE;

endmodule

