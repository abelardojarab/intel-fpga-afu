// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// Frequency monitor for 8 input signals.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_fmon8 #(
    parameter SIM_HURRY = 1'b0,
    parameter SIM_EMULATE = 1'b0
) (
	input clk, 
	input [7:0] din,
	input [2:0] din_sel,
	output [15:0] dout,
	output dout_fresh
);

////////////////////////////
// divide down and cross domain

wire [7:0] prescale;
wire [7:0] prescale_s;

genvar i;
generate
    for (i=0; i<8; i=i+1) begin : lp0
        wire [5:0] local_cnt;
        alt_e100s10_cnt6 ct0 (
            .clk(din[i]),
            .dout(local_cnt)
        );
        defparam ct0 .SIM_EMULATE = SIM_EMULATE;

        assign prescale[i] = local_cnt[5];
        alt_e100s10_sync1r1 sn0 (
            .din_clk(din[i]),
            .din(prescale[i]),
            .dout_clk(clk),
            .dout(prescale_s[i])
        );
        defparam sn0 .SIM_EMULATE = SIM_EMULATE;

    end
endgenerate

////////////////////////////
// select signal to watch

wire sel_prescale;
alt_e100s10_mux8w1t2s1 mx0 (
    .clk(clk),
    .din(prescale_s),
    .sel(din_sel),
    .dout(sel_prescale)
);
defparam mx0 .SIM_EMULATE = SIM_EMULATE;

reg last_sel_prescale = 1'b0;
always @(posedge clk) last_sel_prescale <= sel_prescale;

reg ping = 1'b0;
always @(posedge clk) ping <= sel_prescale ^ last_sel_prescale;

////////////////////////////
// count selected signal

wire sclr;
alt_e100s10_ripple16 rp0 (
    .clk(clk),
    .sclr(sclr),
    .inc(ping),
    .dout(dout)
);
defparam rp0 .SIM_EMULATE = SIM_EMULATE;

////////////////////////////
// regular measuring interval

generate
    if (SIM_HURRY) begin
        // times 100 KHz
        alt_e100s10_metronome32000 mt0 (
            .clk(clk),
            .sclr(1'b0),
            .dout(sclr)
        );
        defparam mt0 .SIM_EMULATE = SIM_EMULATE;

    end
    else begin
        // times 10 KHz
        alt_e100s10_metronome320000 mt0 (
            .clk(clk),
            .sclr(1'b0),
            .dout(sclr)
        );
        defparam mt0 .SIM_EMULATE = SIM_EMULATE;

    end
endgenerate

assign dout_fresh = sclr;
endmodule

