// (C) 2001-2018 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.




`timescale 1ps/1ps

// DESCRIPTION
// MLAB with 16 bit words.  1 addr lines.
// Generated by one of Gregg's toys.   Share And Enjoy.

module alt_e100s10_mlab16a1r1w1 #(
    parameter SIM_EMULATE = 1'b0
) (
    input wclk,
    input [0:0] waddr,
    input [15:0] din,
    input rclk,
    input [0:0] raddr,
    output [15:0] dout
);

////////////////////////////
// handle data bits 15..0

reg [0:0] waddr_m0 = 1'b0 /* synthesis preserve_syn_only */;
always @(posedge wclk) waddr_m0 <= waddr;

reg [15:0] wdata_m0 = 16'b0 /* synthesis preserve_syn_only */;
always @(posedge wclk) wdata_m0 <= din[15:0];

reg [0:0] raddr_m0 = 1'b0 /* synthesis preserve_syn_only */;
always @(posedge rclk) raddr_m0 <= raddr;

alt_e100s10_mlab m0 (
	.wclk(wclk),
	.wena(1'b1),
	.waddr_reg(waddr_m0),
	.wdata_reg(wdata_m0),
	.raddr(raddr_m0),
	.rdata(dout[15:0])
);
defparam m0 .WIDTH = 16;
defparam m0 .ADDR_WIDTH = 1;
defparam m0 .SIM_EMULATE = SIM_EMULATE;

endmodule

